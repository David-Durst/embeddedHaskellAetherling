// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  output [31:0] O_0,
  output [31:0] O_1
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x241_TREADY(dontcare), // @[:@1298.4]
    .io_in_x241_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x241_TID(8'h0),
    .io_in_x241_TDEST(8'h0),
    .io_in_x242_TVALID(valid_down), // @[:@1298.4]
    .io_in_x242_TDATA({O_0,O_1}), // @[:@1298.4]
    .io_in_x242_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x249_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(reset), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule


// End boilerplate
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh27); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh27); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x243_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x518_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x443_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x244_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x245_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x249_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x267_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x492_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x255_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x267_inr_Foreach_kernelx267_inr_Foreach_concrete1( // @[:@5106.2]
  input         clock, // @[:@5107.4]
  input         reset, // @[:@5108.4]
  output        io_in_x245_fifoinpacked_0_wPort_0_en_0, // @[:@5109.4]
  input         io_in_x245_fifoinpacked_0_full, // @[:@5109.4]
  output        io_in_x245_fifoinpacked_0_active_0_in, // @[:@5109.4]
  input         io_in_x245_fifoinpacked_0_active_0_out, // @[:@5109.4]
  input         io_sigsIn_backpressure, // @[:@5109.4]
  input         io_sigsIn_datapathEn, // @[:@5109.4]
  input         io_sigsIn_break, // @[:@5109.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@5109.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5109.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5109.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@5109.4]
  input         io_rr // @[:@5109.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@5143.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@5143.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@5155.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@5155.4]
  wire  x492_sub_1_clock; // @[Math.scala 191:24:@5182.4]
  wire  x492_sub_1_reset; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x492_sub_1_io_a; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x492_sub_1_io_b; // @[Math.scala 191:24:@5182.4]
  wire  x492_sub_1_io_flow; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x492_sub_1_io_result; // @[Math.scala 191:24:@5182.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5192.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5192.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5192.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5192.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5192.4]
  wire  x255_sum_1_clock; // @[Math.scala 150:24:@5201.4]
  wire  x255_sum_1_reset; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x255_sum_1_io_a; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x255_sum_1_io_b; // @[Math.scala 150:24:@5201.4]
  wire  x255_sum_1_io_flow; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x255_sum_1_io_result; // @[Math.scala 150:24:@5201.4]
  wire  x256_sum_1_clock; // @[Math.scala 150:24:@5213.4]
  wire  x256_sum_1_reset; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x256_sum_1_io_a; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x256_sum_1_io_b; // @[Math.scala 150:24:@5213.4]
  wire  x256_sum_1_io_flow; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x256_sum_1_io_result; // @[Math.scala 150:24:@5213.4]
  wire  x494_sum_1_clock; // @[Math.scala 150:24:@5228.4]
  wire  x494_sum_1_reset; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x494_sum_1_io_a; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x494_sum_1_io_b; // @[Math.scala 150:24:@5228.4]
  wire  x494_sum_1_io_flow; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x494_sum_1_io_result; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x259_1_io_b; // @[Math.scala 720:24:@5249.4]
  wire [31:0] x259_1_io_result; // @[Math.scala 720:24:@5249.4]
  wire  x260_sum_1_clock; // @[Math.scala 150:24:@5260.4]
  wire  x260_sum_1_reset; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x260_sum_1_io_a; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x260_sum_1_io_b; // @[Math.scala 150:24:@5260.4]
  wire  x260_sum_1_io_flow; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x260_sum_1_io_result; // @[Math.scala 150:24:@5260.4]
  wire  x497_sum_1_clock; // @[Math.scala 150:24:@5275.4]
  wire  x497_sum_1_reset; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x497_sum_1_io_a; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x497_sum_1_io_b; // @[Math.scala 150:24:@5275.4]
  wire  x497_sum_1_io_flow; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x497_sum_1_io_result; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x263_1_io_b; // @[Math.scala 720:24:@5296.4]
  wire [31:0] x263_1_io_result; // @[Math.scala 720:24:@5296.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5331.4]
  wire  _T_327; // @[sm_x267_inr_Foreach.scala 62:18:@5168.4]
  wire  _T_328; // @[sm_x267_inr_Foreach.scala 62:55:@5169.4]
  wire [31:0] b250_number; // @[Math.scala 723:22:@5148.4 Math.scala 724:14:@5149.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@5173.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@5173.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@5178.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@5178.4]
  wire [31:0] x256_sum_number; // @[Math.scala 154:22:@5219.4 Math.scala 155:14:@5220.4]
  wire [33:0] _GEN_2; // @[Math.scala 461:32:@5224.4]
  wire [33:0] _T_353; // @[Math.scala 461:32:@5224.4]
  wire [31:0] x494_sum_number; // @[Math.scala 154:22:@5234.4 Math.scala 155:14:@5235.4]
  wire [31:0] _T_364; // @[Math.scala 406:49:@5241.4]
  wire [31:0] _T_366; // @[Math.scala 406:56:@5243.4]
  wire [31:0] _T_367; // @[Math.scala 406:56:@5244.4]
  wire [31:0] x260_sum_number; // @[Math.scala 154:22:@5266.4 Math.scala 155:14:@5267.4]
  wire [33:0] _GEN_3; // @[Math.scala 461:32:@5271.4]
  wire [33:0] _T_381; // @[Math.scala 461:32:@5271.4]
  wire [31:0] x497_sum_number; // @[Math.scala 154:22:@5281.4 Math.scala 155:14:@5282.4]
  wire [31:0] _T_392; // @[Math.scala 406:49:@5288.4]
  wire [31:0] _T_394; // @[Math.scala 406:56:@5290.4]
  wire [31:0] _T_395; // @[Math.scala 406:56:@5291.4]
  wire  _T_415; // @[sm_x267_inr_Foreach.scala 103:131:@5328.4]
  wire  _T_419; // @[package.scala 96:25:@5336.4 package.scala 96:25:@5337.4]
  wire  _T_421; // @[implicits.scala 55:10:@5338.4]
  wire  _T_422; // @[sm_x267_inr_Foreach.scala 103:148:@5339.4]
  wire  _T_424; // @[sm_x267_inr_Foreach.scala 103:236:@5341.4]
  wire  _T_425; // @[sm_x267_inr_Foreach.scala 103:255:@5342.4]
  wire  x521_b252_D4; // @[package.scala 96:25:@5316.4 package.scala 96:25:@5317.4]
  wire  _T_428; // @[sm_x267_inr_Foreach.scala 103:291:@5344.4]
  wire  x522_b253_D4; // @[package.scala 96:25:@5325.4 package.scala 96:25:@5326.4]
  _ _ ( // @[Math.scala 720:24:@5143.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@5155.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x492_sub x492_sub_1 ( // @[Math.scala 191:24:@5182.4]
    .clock(x492_sub_1_clock),
    .reset(x492_sub_1_reset),
    .io_a(x492_sub_1_io_a),
    .io_b(x492_sub_1_io_b),
    .io_flow(x492_sub_1_io_flow),
    .io_result(x492_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@5192.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x255_sum x255_sum_1 ( // @[Math.scala 150:24:@5201.4]
    .clock(x255_sum_1_clock),
    .reset(x255_sum_1_reset),
    .io_a(x255_sum_1_io_a),
    .io_b(x255_sum_1_io_b),
    .io_flow(x255_sum_1_io_flow),
    .io_result(x255_sum_1_io_result)
  );
  x255_sum x256_sum_1 ( // @[Math.scala 150:24:@5213.4]
    .clock(x256_sum_1_clock),
    .reset(x256_sum_1_reset),
    .io_a(x256_sum_1_io_a),
    .io_b(x256_sum_1_io_b),
    .io_flow(x256_sum_1_io_flow),
    .io_result(x256_sum_1_io_result)
  );
  x255_sum x494_sum_1 ( // @[Math.scala 150:24:@5228.4]
    .clock(x494_sum_1_clock),
    .reset(x494_sum_1_reset),
    .io_a(x494_sum_1_io_a),
    .io_b(x494_sum_1_io_b),
    .io_flow(x494_sum_1_io_flow),
    .io_result(x494_sum_1_io_result)
  );
  _ x259_1 ( // @[Math.scala 720:24:@5249.4]
    .io_b(x259_1_io_b),
    .io_result(x259_1_io_result)
  );
  x255_sum x260_sum_1 ( // @[Math.scala 150:24:@5260.4]
    .clock(x260_sum_1_clock),
    .reset(x260_sum_1_reset),
    .io_a(x260_sum_1_io_a),
    .io_b(x260_sum_1_io_b),
    .io_flow(x260_sum_1_io_flow),
    .io_result(x260_sum_1_io_result)
  );
  x255_sum x497_sum_1 ( // @[Math.scala 150:24:@5275.4]
    .clock(x497_sum_1_clock),
    .reset(x497_sum_1_reset),
    .io_a(x497_sum_1_io_a),
    .io_b(x497_sum_1_io_b),
    .io_flow(x497_sum_1_io_flow),
    .io_result(x497_sum_1_io_result)
  );
  _ x263_1 ( // @[Math.scala 720:24:@5296.4]
    .io_b(x263_1_io_b),
    .io_result(x263_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@5311.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@5320.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@5331.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x245_fifoinpacked_0_full; // @[sm_x267_inr_Foreach.scala 62:18:@5168.4]
  assign _T_328 = ~ io_in_x245_fifoinpacked_0_active_0_out; // @[sm_x267_inr_Foreach.scala 62:55:@5169.4]
  assign b250_number = __io_result; // @[Math.scala 723:22:@5148.4 Math.scala 724:14:@5149.4]
  assign _GEN_0 = {{11'd0}, b250_number}; // @[Math.scala 461:32:@5173.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@5173.4]
  assign _GEN_1 = {{7'd0}, b250_number}; // @[Math.scala 461:32:@5178.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@5178.4]
  assign x256_sum_number = x256_sum_1_io_result; // @[Math.scala 154:22:@5219.4 Math.scala 155:14:@5220.4]
  assign _GEN_2 = {{2'd0}, x256_sum_number}; // @[Math.scala 461:32:@5224.4]
  assign _T_353 = _GEN_2 << 2; // @[Math.scala 461:32:@5224.4]
  assign x494_sum_number = x494_sum_1_io_result; // @[Math.scala 154:22:@5234.4 Math.scala 155:14:@5235.4]
  assign _T_364 = $signed(x494_sum_number); // @[Math.scala 406:49:@5241.4]
  assign _T_366 = $signed(_T_364) & $signed(32'shff); // @[Math.scala 406:56:@5243.4]
  assign _T_367 = $signed(_T_366); // @[Math.scala 406:56:@5244.4]
  assign x260_sum_number = x260_sum_1_io_result; // @[Math.scala 154:22:@5266.4 Math.scala 155:14:@5267.4]
  assign _GEN_3 = {{2'd0}, x260_sum_number}; // @[Math.scala 461:32:@5271.4]
  assign _T_381 = _GEN_3 << 2; // @[Math.scala 461:32:@5271.4]
  assign x497_sum_number = x497_sum_1_io_result; // @[Math.scala 154:22:@5281.4 Math.scala 155:14:@5282.4]
  assign _T_392 = $signed(x497_sum_number); // @[Math.scala 406:49:@5288.4]
  assign _T_394 = $signed(_T_392) & $signed(32'shff); // @[Math.scala 406:56:@5290.4]
  assign _T_395 = $signed(_T_394); // @[Math.scala 406:56:@5291.4]
  assign _T_415 = ~ io_sigsIn_break; // @[sm_x267_inr_Foreach.scala 103:131:@5328.4]
  assign _T_419 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@5336.4 package.scala 96:25:@5337.4]
  assign _T_421 = io_rr ? _T_419 : 1'h0; // @[implicits.scala 55:10:@5338.4]
  assign _T_422 = _T_415 & _T_421; // @[sm_x267_inr_Foreach.scala 103:148:@5339.4]
  assign _T_424 = _T_422 & _T_415; // @[sm_x267_inr_Foreach.scala 103:236:@5341.4]
  assign _T_425 = _T_424 & io_sigsIn_backpressure; // @[sm_x267_inr_Foreach.scala 103:255:@5342.4]
  assign x521_b252_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5316.4 package.scala 96:25:@5317.4]
  assign _T_428 = _T_425 & x521_b252_D4; // @[sm_x267_inr_Foreach.scala 103:291:@5344.4]
  assign x522_b253_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5325.4 package.scala 96:25:@5326.4]
  assign io_in_x245_fifoinpacked_0_wPort_0_en_0 = _T_428 & x522_b253_D4; // @[MemInterfaceType.scala 93:57:@5348.4]
  assign io_in_x245_fifoinpacked_0_active_0_in = x521_b252_D4 & x522_b253_D4; // @[MemInterfaceType.scala 147:18:@5351.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@5146.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@5158.4]
  assign x492_sub_1_clock = clock; // @[:@5183.4]
  assign x492_sub_1_reset = reset; // @[:@5184.4]
  assign x492_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@5185.4]
  assign x492_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@5186.4]
  assign x492_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@5187.4]
  assign RetimeWrapper_clock = clock; // @[:@5193.4]
  assign RetimeWrapper_reset = reset; // @[:@5194.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5196.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@5195.4]
  assign x255_sum_1_clock = clock; // @[:@5202.4]
  assign x255_sum_1_reset = reset; // @[:@5203.4]
  assign x255_sum_1_io_a = x492_sub_1_io_result; // @[Math.scala 151:17:@5204.4]
  assign x255_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@5205.4]
  assign x255_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5206.4]
  assign x256_sum_1_clock = clock; // @[:@5214.4]
  assign x256_sum_1_reset = reset; // @[:@5215.4]
  assign x256_sum_1_io_a = x255_sum_1_io_result; // @[Math.scala 151:17:@5216.4]
  assign x256_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@5217.4]
  assign x256_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5218.4]
  assign x494_sum_1_clock = clock; // @[:@5229.4]
  assign x494_sum_1_reset = reset; // @[:@5230.4]
  assign x494_sum_1_io_a = _T_353[31:0]; // @[Math.scala 151:17:@5231.4]
  assign x494_sum_1_io_b = x256_sum_1_io_result; // @[Math.scala 152:17:@5232.4]
  assign x494_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5233.4]
  assign x259_1_io_b = $unsigned(_T_367); // @[Math.scala 721:17:@5252.4]
  assign x260_sum_1_clock = clock; // @[:@5261.4]
  assign x260_sum_1_reset = reset; // @[:@5262.4]
  assign x260_sum_1_io_a = x255_sum_1_io_result; // @[Math.scala 151:17:@5263.4]
  assign x260_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@5264.4]
  assign x260_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5265.4]
  assign x497_sum_1_clock = clock; // @[:@5276.4]
  assign x497_sum_1_reset = reset; // @[:@5277.4]
  assign x497_sum_1_io_a = _T_381[31:0]; // @[Math.scala 151:17:@5278.4]
  assign x497_sum_1_io_b = x260_sum_1_io_result; // @[Math.scala 152:17:@5279.4]
  assign x497_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5280.4]
  assign x263_1_io_b = $unsigned(_T_395); // @[Math.scala 721:17:@5299.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5312.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5313.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5315.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@5314.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5321.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5322.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5324.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@5323.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5332.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5333.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5335.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5334.4]
endmodule
module RetimeWrapper_44( // @[:@6469.2]
  input   clock, // @[:@6470.4]
  input   reset, // @[:@6471.4]
  input   io_flow, // @[:@6472.4]
  input   io_in, // @[:@6472.4]
  output  io_out // @[:@6472.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@6474.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6487.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6486.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6485.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6484.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6483.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6481.4]
endmodule
module RetimeWrapper_48( // @[:@6597.2]
  input   clock, // @[:@6598.4]
  input   reset, // @[:@6599.4]
  input   io_flow, // @[:@6600.4]
  input   io_in, // @[:@6600.4]
  output  io_out // @[:@6600.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(39)) sr ( // @[RetimeShiftRegister.scala 15:20:@6602.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6615.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6614.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6613.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6612.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6611.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6609.4]
endmodule
module x441_inr_Foreach_SAMPLER_BOX_sm( // @[:@6617.2]
  input   clock, // @[:@6618.4]
  input   reset, // @[:@6619.4]
  input   io_enable, // @[:@6620.4]
  output  io_done, // @[:@6620.4]
  output  io_doneLatch, // @[:@6620.4]
  input   io_ctrDone, // @[:@6620.4]
  output  io_datapathEn, // @[:@6620.4]
  output  io_ctrInc, // @[:@6620.4]
  output  io_ctrRst, // @[:@6620.4]
  input   io_parentAck, // @[:@6620.4]
  input   io_backpressure, // @[:@6620.4]
  input   io_break // @[:@6620.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6622.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6622.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6625.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6625.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6717.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6630.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6631.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6632.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6633.4]
  wire  _T_100; // @[package.scala 100:49:@6650.4]
  reg  _T_103; // @[package.scala 48:56:@6651.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6664.4 package.scala 96:25:@6665.4]
  wire  _T_110; // @[package.scala 100:49:@6666.4]
  reg  _T_113; // @[package.scala 48:56:@6667.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6669.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6674.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6675.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6678.4]
  wire  _T_124; // @[package.scala 96:25:@6686.4 package.scala 96:25:@6687.4]
  wire  _T_126; // @[package.scala 100:49:@6688.4]
  reg  _T_129; // @[package.scala 48:56:@6689.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6711.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6713.4]
  reg  _T_153; // @[package.scala 48:56:@6714.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6722.4 package.scala 96:25:@6723.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6724.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6725.4]
  SRFF active ( // @[Controllers.scala 261:22:@6622.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6625.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@6659.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_1 ( // @[package.scala 93:22:@6681.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6693.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6701.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_4 ( // @[package.scala 93:22:@6717.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6630.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6631.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6632.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6633.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6650.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6664.4 package.scala 96:25:@6665.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6666.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6669.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6674.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6675.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6678.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6686.4 package.scala 96:25:@6687.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6688.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6713.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6722.4 package.scala 96:25:@6723.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6724.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6725.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6692.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6727.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6677.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6680.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6672.4]
  assign active_clock = clock; // @[:@6623.4]
  assign active_reset = reset; // @[:@6624.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6635.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6639.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6640.4]
  assign done_clock = clock; // @[:@6626.4]
  assign done_reset = reset; // @[:@6627.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6655.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6648.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6649.4]
  assign RetimeWrapper_clock = clock; // @[:@6660.4]
  assign RetimeWrapper_reset = reset; // @[:@6661.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6663.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6662.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6682.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6683.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6685.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6684.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6694.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6695.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6697.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6696.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6702.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6703.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6705.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6704.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6718.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6719.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6721.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6720.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_52( // @[:@6918.2]
  input         clock, // @[:@6919.4]
  input         reset, // @[:@6920.4]
  input         io_flow, // @[:@6921.4]
  input  [63:0] io_in, // @[:@6921.4]
  output [63:0] io_out // @[:@6921.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6923.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6936.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6935.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@6934.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6933.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6932.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6930.4]
endmodule
module SRAM_1( // @[:@6954.2]
  input         clock, // @[:@6955.4]
  input         reset, // @[:@6956.4]
  input  [8:0]  io_raddr, // @[:@6957.4]
  input         io_wen, // @[:@6957.4]
  input  [8:0]  io_waddr, // @[:@6957.4]
  input  [31:0] io_wdata, // @[:@6957.4]
  output [31:0] io_rdata, // @[:@6957.4]
  input         io_backpressure // @[:@6957.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6959.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6959.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6959.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6959.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6977.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6978.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6979.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6981.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(480), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6959.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6977.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6978.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6986.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6973.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6974.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6971.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6976.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6975.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6972.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6970.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6969.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_53( // @[:@7000.2]
  input        clock, // @[:@7001.4]
  input        reset, // @[:@7002.4]
  input        io_flow, // @[:@7003.4]
  input  [8:0] io_in, // @[:@7003.4]
  output [8:0] io_out // @[:@7003.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7005.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7018.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7017.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@7016.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7015.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7014.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7012.4]
endmodule
module Mem1D_5( // @[:@7020.2]
  input         clock, // @[:@7021.4]
  input         reset, // @[:@7022.4]
  input  [8:0]  io_r_ofs_0, // @[:@7023.4]
  input         io_r_backpressure, // @[:@7023.4]
  input  [8:0]  io_w_ofs_0, // @[:@7023.4]
  input  [31:0] io_w_data_0, // @[:@7023.4]
  input         io_w_en_0, // @[:@7023.4]
  output [31:0] io_output // @[:@7023.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7030.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7030.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7030.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7030.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7030.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@7025.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@7027.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_53 RetimeWrapper ( // @[package.scala 93:22:@7030.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h1e0; // @[MemPrimitives.scala 702:32:@7025.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@7043.4]
  assign SRAM_clock = clock; // @[:@7028.4]
  assign SRAM_reset = reset; // @[:@7029.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@7037.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@7040.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@7038.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@7041.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@7042.4]
  assign RetimeWrapper_clock = clock; // @[:@7031.4]
  assign RetimeWrapper_reset = reset; // @[:@7032.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@7034.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@7033.4]
endmodule
module StickySelects_1( // @[:@8650.2]
  input   clock, // @[:@8651.4]
  input   reset, // @[:@8652.4]
  input   io_ins_0, // @[:@8653.4]
  input   io_ins_1, // @[:@8653.4]
  input   io_ins_2, // @[:@8653.4]
  input   io_ins_3, // @[:@8653.4]
  input   io_ins_4, // @[:@8653.4]
  input   io_ins_5, // @[:@8653.4]
  output  io_outs_0, // @[:@8653.4]
  output  io_outs_1, // @[:@8653.4]
  output  io_outs_2, // @[:@8653.4]
  output  io_outs_3, // @[:@8653.4]
  output  io_outs_4, // @[:@8653.4]
  output  io_outs_5 // @[:@8653.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@8655.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@8656.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@8657.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@8658.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@8659.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@8660.4]
  reg [31:0] _RAND_5;
  wire  _T_35; // @[StickySelects.scala 47:46:@8661.4]
  wire  _T_36; // @[StickySelects.scala 47:46:@8662.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@8663.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@8664.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@8665.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@8666.4]
  wire  _T_41; // @[StickySelects.scala 47:46:@8668.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@8669.4]
  wire  _T_43; // @[StickySelects.scala 47:46:@8670.4]
  wire  _T_44; // @[StickySelects.scala 47:46:@8671.4]
  wire  _T_45; // @[StickySelects.scala 49:53:@8672.4]
  wire  _T_46; // @[StickySelects.scala 49:21:@8673.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@8675.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@8676.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@8677.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@8678.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@8679.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@8680.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@8683.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@8684.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@8685.4]
  wire  _T_57; // @[StickySelects.scala 49:53:@8686.4]
  wire  _T_58; // @[StickySelects.scala 49:21:@8687.4]
  wire  _T_61; // @[StickySelects.scala 47:46:@8691.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@8692.4]
  wire  _T_63; // @[StickySelects.scala 49:53:@8693.4]
  wire  _T_64; // @[StickySelects.scala 49:21:@8694.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@8699.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@8700.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@8701.4]
  assign _T_35 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@8661.4]
  assign _T_36 = _T_35 | io_ins_3; // @[StickySelects.scala 47:46:@8662.4]
  assign _T_37 = _T_36 | io_ins_4; // @[StickySelects.scala 47:46:@8663.4]
  assign _T_38 = _T_37 | io_ins_5; // @[StickySelects.scala 47:46:@8664.4]
  assign _T_39 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@8665.4]
  assign _T_40 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 49:21:@8666.4]
  assign _T_41 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@8668.4]
  assign _T_42 = _T_41 | io_ins_3; // @[StickySelects.scala 47:46:@8669.4]
  assign _T_43 = _T_42 | io_ins_4; // @[StickySelects.scala 47:46:@8670.4]
  assign _T_44 = _T_43 | io_ins_5; // @[StickySelects.scala 47:46:@8671.4]
  assign _T_45 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@8672.4]
  assign _T_46 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 49:21:@8673.4]
  assign _T_47 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@8675.4]
  assign _T_48 = _T_47 | io_ins_3; // @[StickySelects.scala 47:46:@8676.4]
  assign _T_49 = _T_48 | io_ins_4; // @[StickySelects.scala 47:46:@8677.4]
  assign _T_50 = _T_49 | io_ins_5; // @[StickySelects.scala 47:46:@8678.4]
  assign _T_51 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@8679.4]
  assign _T_52 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 49:21:@8680.4]
  assign _T_54 = _T_47 | io_ins_2; // @[StickySelects.scala 47:46:@8683.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@8684.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@8685.4]
  assign _T_57 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@8686.4]
  assign _T_58 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 49:21:@8687.4]
  assign _T_61 = _T_54 | io_ins_3; // @[StickySelects.scala 47:46:@8691.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 47:46:@8692.4]
  assign _T_63 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@8693.4]
  assign _T_64 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 49:21:@8694.4]
  assign _T_68 = _T_61 | io_ins_4; // @[StickySelects.scala 47:46:@8699.4]
  assign _T_69 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@8700.4]
  assign _T_70 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 49:21:@8701.4]
  assign io_outs_0 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 53:57:@8703.4]
  assign io_outs_1 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 53:57:@8704.4]
  assign io_outs_2 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 53:57:@8705.4]
  assign io_outs_3 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 53:57:@8706.4]
  assign io_outs_4 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 53:57:@8707.4]
  assign io_outs_5 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 53:57:@8708.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_39;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_45;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_51;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_56) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_57;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_62) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_63;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_69;
      end
    end
  end
endmodule
module x278_lb_0( // @[:@12682.2]
  input         clock, // @[:@12683.4]
  input         reset, // @[:@12684.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@12685.4]
  input         io_rPort_11_en_0, // @[:@12685.4]
  input         io_rPort_11_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_11_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@12685.4]
  input         io_rPort_10_en_0, // @[:@12685.4]
  input         io_rPort_10_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_10_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@12685.4]
  input         io_rPort_9_en_0, // @[:@12685.4]
  input         io_rPort_9_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_9_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@12685.4]
  input         io_rPort_8_en_0, // @[:@12685.4]
  input         io_rPort_8_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_8_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@12685.4]
  input         io_rPort_7_en_0, // @[:@12685.4]
  input         io_rPort_7_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_7_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@12685.4]
  input         io_rPort_6_en_0, // @[:@12685.4]
  input         io_rPort_6_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_6_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@12685.4]
  input         io_rPort_5_en_0, // @[:@12685.4]
  input         io_rPort_5_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_5_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@12685.4]
  input         io_rPort_4_en_0, // @[:@12685.4]
  input         io_rPort_4_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_4_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@12685.4]
  input         io_rPort_3_en_0, // @[:@12685.4]
  input         io_rPort_3_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_3_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@12685.4]
  input         io_rPort_2_en_0, // @[:@12685.4]
  input         io_rPort_2_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_2_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@12685.4]
  input         io_rPort_1_en_0, // @[:@12685.4]
  input         io_rPort_1_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_1_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@12685.4]
  input         io_rPort_0_en_0, // @[:@12685.4]
  input         io_rPort_0_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_0_output_0, // @[:@12685.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@12685.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@12685.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@12685.4]
  input  [31:0] io_wPort_1_data_0, // @[:@12685.4]
  input         io_wPort_1_en_0, // @[:@12685.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@12685.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12685.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@12685.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12685.4]
  input         io_wPort_0_en_0 // @[:@12685.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15353.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@13032.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@13033.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@13034.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@13035.4]
  wire [41:0] _T_450; // @[Cat.scala 30:58:@13037.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@13044.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@13045.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@13046.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@13047.4]
  wire [41:0] _T_461; // @[Cat.scala 30:58:@13049.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@13057.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@13058.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@13059.4]
  wire [41:0] _T_472; // @[Cat.scala 30:58:@13061.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@13069.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@13070.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@13071.4]
  wire [41:0] _T_483; // @[Cat.scala 30:58:@13073.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@13080.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@13082.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@13083.4]
  wire [41:0] _T_494; // @[Cat.scala 30:58:@13085.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@13092.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@13094.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@13095.4]
  wire [41:0] _T_505; // @[Cat.scala 30:58:@13097.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@13106.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@13107.4]
  wire [41:0] _T_516; // @[Cat.scala 30:58:@13109.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@13118.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@13119.4]
  wire [41:0] _T_527; // @[Cat.scala 30:58:@13121.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@13128.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@13130.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@13131.4]
  wire [41:0] _T_538; // @[Cat.scala 30:58:@13133.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@13140.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@13142.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@13143.4]
  wire [41:0] _T_549; // @[Cat.scala 30:58:@13145.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@13154.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@13155.4]
  wire [41:0] _T_560; // @[Cat.scala 30:58:@13157.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@13166.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@13167.4]
  wire [41:0] _T_571; // @[Cat.scala 30:58:@13169.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@13176.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@13178.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@13179.4]
  wire [41:0] _T_582; // @[Cat.scala 30:58:@13181.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@13188.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@13190.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@13191.4]
  wire [41:0] _T_593; // @[Cat.scala 30:58:@13193.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@13202.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@13203.4]
  wire [41:0] _T_604; // @[Cat.scala 30:58:@13205.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@13214.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@13215.4]
  wire [41:0] _T_615; // @[Cat.scala 30:58:@13217.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@13224.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@13225.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@13226.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@13228.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@13229.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@13230.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@13232.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@13233.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@13234.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@13236.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13237.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@13238.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@13240.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13241.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13242.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@13244.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13245.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13246.4]
  wire  _T_655; // @[MemPrimitives.scala 126:35:@13257.4]
  wire  _T_656; // @[MemPrimitives.scala 126:35:@13258.4]
  wire  _T_657; // @[MemPrimitives.scala 126:35:@13259.4]
  wire  _T_658; // @[MemPrimitives.scala 126:35:@13260.4]
  wire  _T_659; // @[MemPrimitives.scala 126:35:@13261.4]
  wire  _T_660; // @[MemPrimitives.scala 126:35:@13262.4]
  wire [10:0] _T_662; // @[Cat.scala 30:58:@13264.4]
  wire [10:0] _T_664; // @[Cat.scala 30:58:@13266.4]
  wire [10:0] _T_666; // @[Cat.scala 30:58:@13268.4]
  wire [10:0] _T_668; // @[Cat.scala 30:58:@13270.4]
  wire [10:0] _T_670; // @[Cat.scala 30:58:@13272.4]
  wire [10:0] _T_672; // @[Cat.scala 30:58:@13274.4]
  wire [10:0] _T_673; // @[Mux.scala 31:69:@13275.4]
  wire [10:0] _T_674; // @[Mux.scala 31:69:@13276.4]
  wire [10:0] _T_675; // @[Mux.scala 31:69:@13277.4]
  wire [10:0] _T_676; // @[Mux.scala 31:69:@13278.4]
  wire [10:0] _T_677; // @[Mux.scala 31:69:@13279.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13286.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@13287.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@13290.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@13291.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@13294.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@13295.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@13296.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@13298.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@13299.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@13300.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@13302.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@13303.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@13304.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@13306.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@13307.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@13308.4]
  wire  _T_717; // @[MemPrimitives.scala 126:35:@13319.4]
  wire  _T_718; // @[MemPrimitives.scala 126:35:@13320.4]
  wire  _T_719; // @[MemPrimitives.scala 126:35:@13321.4]
  wire  _T_720; // @[MemPrimitives.scala 126:35:@13322.4]
  wire  _T_721; // @[MemPrimitives.scala 126:35:@13323.4]
  wire  _T_722; // @[MemPrimitives.scala 126:35:@13324.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@13326.4]
  wire [10:0] _T_726; // @[Cat.scala 30:58:@13328.4]
  wire [10:0] _T_728; // @[Cat.scala 30:58:@13330.4]
  wire [10:0] _T_730; // @[Cat.scala 30:58:@13332.4]
  wire [10:0] _T_732; // @[Cat.scala 30:58:@13334.4]
  wire [10:0] _T_734; // @[Cat.scala 30:58:@13336.4]
  wire [10:0] _T_735; // @[Mux.scala 31:69:@13337.4]
  wire [10:0] _T_736; // @[Mux.scala 31:69:@13338.4]
  wire [10:0] _T_737; // @[Mux.scala 31:69:@13339.4]
  wire [10:0] _T_738; // @[Mux.scala 31:69:@13340.4]
  wire [10:0] _T_739; // @[Mux.scala 31:69:@13341.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@13349.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@13350.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@13353.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@13354.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@13357.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@13358.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@13361.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@13362.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@13365.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@13366.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@13369.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@13370.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@13381.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@13382.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@13383.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@13384.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@13385.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@13386.4]
  wire [10:0] _T_786; // @[Cat.scala 30:58:@13388.4]
  wire [10:0] _T_788; // @[Cat.scala 30:58:@13390.4]
  wire [10:0] _T_790; // @[Cat.scala 30:58:@13392.4]
  wire [10:0] _T_792; // @[Cat.scala 30:58:@13394.4]
  wire [10:0] _T_794; // @[Cat.scala 30:58:@13396.4]
  wire [10:0] _T_796; // @[Cat.scala 30:58:@13398.4]
  wire [10:0] _T_797; // @[Mux.scala 31:69:@13399.4]
  wire [10:0] _T_798; // @[Mux.scala 31:69:@13400.4]
  wire [10:0] _T_799; // @[Mux.scala 31:69:@13401.4]
  wire [10:0] _T_800; // @[Mux.scala 31:69:@13402.4]
  wire [10:0] _T_801; // @[Mux.scala 31:69:@13403.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@13411.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@13412.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@13415.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@13416.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@13419.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@13420.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@13423.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@13424.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@13427.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@13428.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@13431.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@13432.4]
  wire  _T_841; // @[MemPrimitives.scala 126:35:@13443.4]
  wire  _T_842; // @[MemPrimitives.scala 126:35:@13444.4]
  wire  _T_843; // @[MemPrimitives.scala 126:35:@13445.4]
  wire  _T_844; // @[MemPrimitives.scala 126:35:@13446.4]
  wire  _T_845; // @[MemPrimitives.scala 126:35:@13447.4]
  wire  _T_846; // @[MemPrimitives.scala 126:35:@13448.4]
  wire [10:0] _T_848; // @[Cat.scala 30:58:@13450.4]
  wire [10:0] _T_850; // @[Cat.scala 30:58:@13452.4]
  wire [10:0] _T_852; // @[Cat.scala 30:58:@13454.4]
  wire [10:0] _T_854; // @[Cat.scala 30:58:@13456.4]
  wire [10:0] _T_856; // @[Cat.scala 30:58:@13458.4]
  wire [10:0] _T_858; // @[Cat.scala 30:58:@13460.4]
  wire [10:0] _T_859; // @[Mux.scala 31:69:@13461.4]
  wire [10:0] _T_860; // @[Mux.scala 31:69:@13462.4]
  wire [10:0] _T_861; // @[Mux.scala 31:69:@13463.4]
  wire [10:0] _T_862; // @[Mux.scala 31:69:@13464.4]
  wire [10:0] _T_863; // @[Mux.scala 31:69:@13465.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@13472.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@13474.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@13476.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@13478.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@13480.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@13482.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@13484.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@13486.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@13488.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@13490.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@13492.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@13494.4]
  wire  _T_903; // @[MemPrimitives.scala 126:35:@13505.4]
  wire  _T_904; // @[MemPrimitives.scala 126:35:@13506.4]
  wire  _T_905; // @[MemPrimitives.scala 126:35:@13507.4]
  wire  _T_906; // @[MemPrimitives.scala 126:35:@13508.4]
  wire  _T_907; // @[MemPrimitives.scala 126:35:@13509.4]
  wire  _T_908; // @[MemPrimitives.scala 126:35:@13510.4]
  wire [10:0] _T_910; // @[Cat.scala 30:58:@13512.4]
  wire [10:0] _T_912; // @[Cat.scala 30:58:@13514.4]
  wire [10:0] _T_914; // @[Cat.scala 30:58:@13516.4]
  wire [10:0] _T_916; // @[Cat.scala 30:58:@13518.4]
  wire [10:0] _T_918; // @[Cat.scala 30:58:@13520.4]
  wire [10:0] _T_920; // @[Cat.scala 30:58:@13522.4]
  wire [10:0] _T_921; // @[Mux.scala 31:69:@13523.4]
  wire [10:0] _T_922; // @[Mux.scala 31:69:@13524.4]
  wire [10:0] _T_923; // @[Mux.scala 31:69:@13525.4]
  wire [10:0] _T_924; // @[Mux.scala 31:69:@13526.4]
  wire [10:0] _T_925; // @[Mux.scala 31:69:@13527.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@13534.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@13536.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@13538.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@13540.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@13542.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@13544.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@13546.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@13548.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@13550.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@13552.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@13554.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@13556.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13567.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13568.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13569.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13570.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13571.4]
  wire  _T_970; // @[MemPrimitives.scala 126:35:@13572.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@13574.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@13576.4]
  wire [10:0] _T_976; // @[Cat.scala 30:58:@13578.4]
  wire [10:0] _T_978; // @[Cat.scala 30:58:@13580.4]
  wire [10:0] _T_980; // @[Cat.scala 30:58:@13582.4]
  wire [10:0] _T_982; // @[Cat.scala 30:58:@13584.4]
  wire [10:0] _T_983; // @[Mux.scala 31:69:@13585.4]
  wire [10:0] _T_984; // @[Mux.scala 31:69:@13586.4]
  wire [10:0] _T_985; // @[Mux.scala 31:69:@13587.4]
  wire [10:0] _T_986; // @[Mux.scala 31:69:@13588.4]
  wire [10:0] _T_987; // @[Mux.scala 31:69:@13589.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@13598.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@13602.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@13606.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@13610.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@13614.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@13618.4]
  wire  _T_1027; // @[MemPrimitives.scala 126:35:@13629.4]
  wire  _T_1028; // @[MemPrimitives.scala 126:35:@13630.4]
  wire  _T_1029; // @[MemPrimitives.scala 126:35:@13631.4]
  wire  _T_1030; // @[MemPrimitives.scala 126:35:@13632.4]
  wire  _T_1031; // @[MemPrimitives.scala 126:35:@13633.4]
  wire  _T_1032; // @[MemPrimitives.scala 126:35:@13634.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@13636.4]
  wire [10:0] _T_1036; // @[Cat.scala 30:58:@13638.4]
  wire [10:0] _T_1038; // @[Cat.scala 30:58:@13640.4]
  wire [10:0] _T_1040; // @[Cat.scala 30:58:@13642.4]
  wire [10:0] _T_1042; // @[Cat.scala 30:58:@13644.4]
  wire [10:0] _T_1044; // @[Cat.scala 30:58:@13646.4]
  wire [10:0] _T_1045; // @[Mux.scala 31:69:@13647.4]
  wire [10:0] _T_1046; // @[Mux.scala 31:69:@13648.4]
  wire [10:0] _T_1047; // @[Mux.scala 31:69:@13649.4]
  wire [10:0] _T_1048; // @[Mux.scala 31:69:@13650.4]
  wire [10:0] _T_1049; // @[Mux.scala 31:69:@13651.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@13660.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@13664.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@13668.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@13672.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@13676.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@13680.4]
  wire  _T_1089; // @[MemPrimitives.scala 126:35:@13691.4]
  wire  _T_1090; // @[MemPrimitives.scala 126:35:@13692.4]
  wire  _T_1091; // @[MemPrimitives.scala 126:35:@13693.4]
  wire  _T_1092; // @[MemPrimitives.scala 126:35:@13694.4]
  wire  _T_1093; // @[MemPrimitives.scala 126:35:@13695.4]
  wire  _T_1094; // @[MemPrimitives.scala 126:35:@13696.4]
  wire [10:0] _T_1096; // @[Cat.scala 30:58:@13698.4]
  wire [10:0] _T_1098; // @[Cat.scala 30:58:@13700.4]
  wire [10:0] _T_1100; // @[Cat.scala 30:58:@13702.4]
  wire [10:0] _T_1102; // @[Cat.scala 30:58:@13704.4]
  wire [10:0] _T_1104; // @[Cat.scala 30:58:@13706.4]
  wire [10:0] _T_1106; // @[Cat.scala 30:58:@13708.4]
  wire [10:0] _T_1107; // @[Mux.scala 31:69:@13709.4]
  wire [10:0] _T_1108; // @[Mux.scala 31:69:@13710.4]
  wire [10:0] _T_1109; // @[Mux.scala 31:69:@13711.4]
  wire [10:0] _T_1110; // @[Mux.scala 31:69:@13712.4]
  wire [10:0] _T_1111; // @[Mux.scala 31:69:@13713.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@13720.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13722.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@13724.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13726.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@13728.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13730.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@13732.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13734.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@13736.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13738.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@13740.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@13742.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13753.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13754.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13755.4]
  wire  _T_1154; // @[MemPrimitives.scala 126:35:@13756.4]
  wire  _T_1155; // @[MemPrimitives.scala 126:35:@13757.4]
  wire  _T_1156; // @[MemPrimitives.scala 126:35:@13758.4]
  wire [10:0] _T_1158; // @[Cat.scala 30:58:@13760.4]
  wire [10:0] _T_1160; // @[Cat.scala 30:58:@13762.4]
  wire [10:0] _T_1162; // @[Cat.scala 30:58:@13764.4]
  wire [10:0] _T_1164; // @[Cat.scala 30:58:@13766.4]
  wire [10:0] _T_1166; // @[Cat.scala 30:58:@13768.4]
  wire [10:0] _T_1168; // @[Cat.scala 30:58:@13770.4]
  wire [10:0] _T_1169; // @[Mux.scala 31:69:@13771.4]
  wire [10:0] _T_1170; // @[Mux.scala 31:69:@13772.4]
  wire [10:0] _T_1171; // @[Mux.scala 31:69:@13773.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@13774.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@13775.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@13782.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@13784.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@13786.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13788.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@13790.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13792.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@13794.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13796.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@13798.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13800.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@13802.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13804.4]
  wire  _T_1213; // @[MemPrimitives.scala 126:35:@13815.4]
  wire  _T_1214; // @[MemPrimitives.scala 126:35:@13816.4]
  wire  _T_1215; // @[MemPrimitives.scala 126:35:@13817.4]
  wire  _T_1216; // @[MemPrimitives.scala 126:35:@13818.4]
  wire  _T_1217; // @[MemPrimitives.scala 126:35:@13819.4]
  wire  _T_1218; // @[MemPrimitives.scala 126:35:@13820.4]
  wire [10:0] _T_1220; // @[Cat.scala 30:58:@13822.4]
  wire [10:0] _T_1222; // @[Cat.scala 30:58:@13824.4]
  wire [10:0] _T_1224; // @[Cat.scala 30:58:@13826.4]
  wire [10:0] _T_1226; // @[Cat.scala 30:58:@13828.4]
  wire [10:0] _T_1228; // @[Cat.scala 30:58:@13830.4]
  wire [10:0] _T_1230; // @[Cat.scala 30:58:@13832.4]
  wire [10:0] _T_1231; // @[Mux.scala 31:69:@13833.4]
  wire [10:0] _T_1232; // @[Mux.scala 31:69:@13834.4]
  wire [10:0] _T_1233; // @[Mux.scala 31:69:@13835.4]
  wire [10:0] _T_1234; // @[Mux.scala 31:69:@13836.4]
  wire [10:0] _T_1235; // @[Mux.scala 31:69:@13837.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@13846.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@13850.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@13854.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@13858.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@13862.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@13866.4]
  wire  _T_1275; // @[MemPrimitives.scala 126:35:@13877.4]
  wire  _T_1276; // @[MemPrimitives.scala 126:35:@13878.4]
  wire  _T_1277; // @[MemPrimitives.scala 126:35:@13879.4]
  wire  _T_1278; // @[MemPrimitives.scala 126:35:@13880.4]
  wire  _T_1279; // @[MemPrimitives.scala 126:35:@13881.4]
  wire  _T_1280; // @[MemPrimitives.scala 126:35:@13882.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@13884.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@13886.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@13888.4]
  wire [10:0] _T_1288; // @[Cat.scala 30:58:@13890.4]
  wire [10:0] _T_1290; // @[Cat.scala 30:58:@13892.4]
  wire [10:0] _T_1292; // @[Cat.scala 30:58:@13894.4]
  wire [10:0] _T_1293; // @[Mux.scala 31:69:@13895.4]
  wire [10:0] _T_1294; // @[Mux.scala 31:69:@13896.4]
  wire [10:0] _T_1295; // @[Mux.scala 31:69:@13897.4]
  wire [10:0] _T_1296; // @[Mux.scala 31:69:@13898.4]
  wire [10:0] _T_1297; // @[Mux.scala 31:69:@13899.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@13908.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@13912.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@13916.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@13920.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@13924.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@13928.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13939.4]
  wire  _T_1338; // @[MemPrimitives.scala 126:35:@13940.4]
  wire  _T_1339; // @[MemPrimitives.scala 126:35:@13941.4]
  wire  _T_1340; // @[MemPrimitives.scala 126:35:@13942.4]
  wire  _T_1341; // @[MemPrimitives.scala 126:35:@13943.4]
  wire  _T_1342; // @[MemPrimitives.scala 126:35:@13944.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@13946.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@13948.4]
  wire [10:0] _T_1348; // @[Cat.scala 30:58:@13950.4]
  wire [10:0] _T_1350; // @[Cat.scala 30:58:@13952.4]
  wire [10:0] _T_1352; // @[Cat.scala 30:58:@13954.4]
  wire [10:0] _T_1354; // @[Cat.scala 30:58:@13956.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@13957.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@13958.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@13959.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@13960.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@13961.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@13968.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@13970.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@13972.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@13974.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@13976.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@13978.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@13980.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@13982.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@13984.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@13986.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@13988.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@13990.4]
  wire  _T_1399; // @[MemPrimitives.scala 126:35:@14001.4]
  wire  _T_1400; // @[MemPrimitives.scala 126:35:@14002.4]
  wire  _T_1401; // @[MemPrimitives.scala 126:35:@14003.4]
  wire  _T_1402; // @[MemPrimitives.scala 126:35:@14004.4]
  wire  _T_1403; // @[MemPrimitives.scala 126:35:@14005.4]
  wire  _T_1404; // @[MemPrimitives.scala 126:35:@14006.4]
  wire [10:0] _T_1406; // @[Cat.scala 30:58:@14008.4]
  wire [10:0] _T_1408; // @[Cat.scala 30:58:@14010.4]
  wire [10:0] _T_1410; // @[Cat.scala 30:58:@14012.4]
  wire [10:0] _T_1412; // @[Cat.scala 30:58:@14014.4]
  wire [10:0] _T_1414; // @[Cat.scala 30:58:@14016.4]
  wire [10:0] _T_1416; // @[Cat.scala 30:58:@14018.4]
  wire [10:0] _T_1417; // @[Mux.scala 31:69:@14019.4]
  wire [10:0] _T_1418; // @[Mux.scala 31:69:@14020.4]
  wire [10:0] _T_1419; // @[Mux.scala 31:69:@14021.4]
  wire [10:0] _T_1420; // @[Mux.scala 31:69:@14022.4]
  wire [10:0] _T_1421; // @[Mux.scala 31:69:@14023.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@14030.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@14032.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@14034.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@14036.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@14038.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@14040.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@14042.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@14044.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@14046.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@14048.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@14050.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@14052.4]
  wire  _T_1461; // @[MemPrimitives.scala 126:35:@14063.4]
  wire  _T_1462; // @[MemPrimitives.scala 126:35:@14064.4]
  wire  _T_1463; // @[MemPrimitives.scala 126:35:@14065.4]
  wire  _T_1464; // @[MemPrimitives.scala 126:35:@14066.4]
  wire  _T_1465; // @[MemPrimitives.scala 126:35:@14067.4]
  wire  _T_1466; // @[MemPrimitives.scala 126:35:@14068.4]
  wire [10:0] _T_1468; // @[Cat.scala 30:58:@14070.4]
  wire [10:0] _T_1470; // @[Cat.scala 30:58:@14072.4]
  wire [10:0] _T_1472; // @[Cat.scala 30:58:@14074.4]
  wire [10:0] _T_1474; // @[Cat.scala 30:58:@14076.4]
  wire [10:0] _T_1476; // @[Cat.scala 30:58:@14078.4]
  wire [10:0] _T_1478; // @[Cat.scala 30:58:@14080.4]
  wire [10:0] _T_1479; // @[Mux.scala 31:69:@14081.4]
  wire [10:0] _T_1480; // @[Mux.scala 31:69:@14082.4]
  wire [10:0] _T_1481; // @[Mux.scala 31:69:@14083.4]
  wire [10:0] _T_1482; // @[Mux.scala 31:69:@14084.4]
  wire [10:0] _T_1483; // @[Mux.scala 31:69:@14085.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@14094.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@14098.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@14102.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@14106.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@14110.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@14114.4]
  wire  _T_1523; // @[MemPrimitives.scala 126:35:@14125.4]
  wire  _T_1524; // @[MemPrimitives.scala 126:35:@14126.4]
  wire  _T_1525; // @[MemPrimitives.scala 126:35:@14127.4]
  wire  _T_1526; // @[MemPrimitives.scala 126:35:@14128.4]
  wire  _T_1527; // @[MemPrimitives.scala 126:35:@14129.4]
  wire  _T_1528; // @[MemPrimitives.scala 126:35:@14130.4]
  wire [10:0] _T_1530; // @[Cat.scala 30:58:@14132.4]
  wire [10:0] _T_1532; // @[Cat.scala 30:58:@14134.4]
  wire [10:0] _T_1534; // @[Cat.scala 30:58:@14136.4]
  wire [10:0] _T_1536; // @[Cat.scala 30:58:@14138.4]
  wire [10:0] _T_1538; // @[Cat.scala 30:58:@14140.4]
  wire [10:0] _T_1540; // @[Cat.scala 30:58:@14142.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@14143.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@14144.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@14145.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@14146.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@14147.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@14156.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@14160.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@14164.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@14168.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@14172.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@14176.4]
  wire  _T_1585; // @[MemPrimitives.scala 126:35:@14187.4]
  wire  _T_1586; // @[MemPrimitives.scala 126:35:@14188.4]
  wire  _T_1587; // @[MemPrimitives.scala 126:35:@14189.4]
  wire  _T_1588; // @[MemPrimitives.scala 126:35:@14190.4]
  wire  _T_1589; // @[MemPrimitives.scala 126:35:@14191.4]
  wire  _T_1590; // @[MemPrimitives.scala 126:35:@14192.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@14194.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@14196.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@14198.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@14200.4]
  wire [10:0] _T_1600; // @[Cat.scala 30:58:@14202.4]
  wire [10:0] _T_1602; // @[Cat.scala 30:58:@14204.4]
  wire [10:0] _T_1603; // @[Mux.scala 31:69:@14205.4]
  wire [10:0] _T_1604; // @[Mux.scala 31:69:@14206.4]
  wire [10:0] _T_1605; // @[Mux.scala 31:69:@14207.4]
  wire [10:0] _T_1606; // @[Mux.scala 31:69:@14208.4]
  wire [10:0] _T_1607; // @[Mux.scala 31:69:@14209.4]
  wire  _T_1671; // @[package.scala 96:25:@14294.4 package.scala 96:25:@14295.4]
  wire [31:0] _T_1675; // @[Mux.scala 31:69:@14304.4]
  wire  _T_1668; // @[package.scala 96:25:@14286.4 package.scala 96:25:@14287.4]
  wire [31:0] _T_1676; // @[Mux.scala 31:69:@14305.4]
  wire  _T_1665; // @[package.scala 96:25:@14278.4 package.scala 96:25:@14279.4]
  wire [31:0] _T_1677; // @[Mux.scala 31:69:@14306.4]
  wire  _T_1662; // @[package.scala 96:25:@14270.4 package.scala 96:25:@14271.4]
  wire [31:0] _T_1678; // @[Mux.scala 31:69:@14307.4]
  wire  _T_1659; // @[package.scala 96:25:@14262.4 package.scala 96:25:@14263.4]
  wire [31:0] _T_1679; // @[Mux.scala 31:69:@14308.4]
  wire  _T_1656; // @[package.scala 96:25:@14254.4 package.scala 96:25:@14255.4]
  wire [31:0] _T_1680; // @[Mux.scala 31:69:@14309.4]
  wire  _T_1653; // @[package.scala 96:25:@14246.4 package.scala 96:25:@14247.4]
  wire  _T_1742; // @[package.scala 96:25:@14390.4 package.scala 96:25:@14391.4]
  wire [31:0] _T_1746; // @[Mux.scala 31:69:@14400.4]
  wire  _T_1739; // @[package.scala 96:25:@14382.4 package.scala 96:25:@14383.4]
  wire [31:0] _T_1747; // @[Mux.scala 31:69:@14401.4]
  wire  _T_1736; // @[package.scala 96:25:@14374.4 package.scala 96:25:@14375.4]
  wire [31:0] _T_1748; // @[Mux.scala 31:69:@14402.4]
  wire  _T_1733; // @[package.scala 96:25:@14366.4 package.scala 96:25:@14367.4]
  wire [31:0] _T_1749; // @[Mux.scala 31:69:@14403.4]
  wire  _T_1730; // @[package.scala 96:25:@14358.4 package.scala 96:25:@14359.4]
  wire [31:0] _T_1750; // @[Mux.scala 31:69:@14404.4]
  wire  _T_1727; // @[package.scala 96:25:@14350.4 package.scala 96:25:@14351.4]
  wire [31:0] _T_1751; // @[Mux.scala 31:69:@14405.4]
  wire  _T_1724; // @[package.scala 96:25:@14342.4 package.scala 96:25:@14343.4]
  wire  _T_1813; // @[package.scala 96:25:@14486.4 package.scala 96:25:@14487.4]
  wire [31:0] _T_1817; // @[Mux.scala 31:69:@14496.4]
  wire  _T_1810; // @[package.scala 96:25:@14478.4 package.scala 96:25:@14479.4]
  wire [31:0] _T_1818; // @[Mux.scala 31:69:@14497.4]
  wire  _T_1807; // @[package.scala 96:25:@14470.4 package.scala 96:25:@14471.4]
  wire [31:0] _T_1819; // @[Mux.scala 31:69:@14498.4]
  wire  _T_1804; // @[package.scala 96:25:@14462.4 package.scala 96:25:@14463.4]
  wire [31:0] _T_1820; // @[Mux.scala 31:69:@14499.4]
  wire  _T_1801; // @[package.scala 96:25:@14454.4 package.scala 96:25:@14455.4]
  wire [31:0] _T_1821; // @[Mux.scala 31:69:@14500.4]
  wire  _T_1798; // @[package.scala 96:25:@14446.4 package.scala 96:25:@14447.4]
  wire [31:0] _T_1822; // @[Mux.scala 31:69:@14501.4]
  wire  _T_1795; // @[package.scala 96:25:@14438.4 package.scala 96:25:@14439.4]
  wire  _T_1884; // @[package.scala 96:25:@14582.4 package.scala 96:25:@14583.4]
  wire [31:0] _T_1888; // @[Mux.scala 31:69:@14592.4]
  wire  _T_1881; // @[package.scala 96:25:@14574.4 package.scala 96:25:@14575.4]
  wire [31:0] _T_1889; // @[Mux.scala 31:69:@14593.4]
  wire  _T_1878; // @[package.scala 96:25:@14566.4 package.scala 96:25:@14567.4]
  wire [31:0] _T_1890; // @[Mux.scala 31:69:@14594.4]
  wire  _T_1875; // @[package.scala 96:25:@14558.4 package.scala 96:25:@14559.4]
  wire [31:0] _T_1891; // @[Mux.scala 31:69:@14595.4]
  wire  _T_1872; // @[package.scala 96:25:@14550.4 package.scala 96:25:@14551.4]
  wire [31:0] _T_1892; // @[Mux.scala 31:69:@14596.4]
  wire  _T_1869; // @[package.scala 96:25:@14542.4 package.scala 96:25:@14543.4]
  wire [31:0] _T_1893; // @[Mux.scala 31:69:@14597.4]
  wire  _T_1866; // @[package.scala 96:25:@14534.4 package.scala 96:25:@14535.4]
  wire  _T_1955; // @[package.scala 96:25:@14678.4 package.scala 96:25:@14679.4]
  wire [31:0] _T_1959; // @[Mux.scala 31:69:@14688.4]
  wire  _T_1952; // @[package.scala 96:25:@14670.4 package.scala 96:25:@14671.4]
  wire [31:0] _T_1960; // @[Mux.scala 31:69:@14689.4]
  wire  _T_1949; // @[package.scala 96:25:@14662.4 package.scala 96:25:@14663.4]
  wire [31:0] _T_1961; // @[Mux.scala 31:69:@14690.4]
  wire  _T_1946; // @[package.scala 96:25:@14654.4 package.scala 96:25:@14655.4]
  wire [31:0] _T_1962; // @[Mux.scala 31:69:@14691.4]
  wire  _T_1943; // @[package.scala 96:25:@14646.4 package.scala 96:25:@14647.4]
  wire [31:0] _T_1963; // @[Mux.scala 31:69:@14692.4]
  wire  _T_1940; // @[package.scala 96:25:@14638.4 package.scala 96:25:@14639.4]
  wire [31:0] _T_1964; // @[Mux.scala 31:69:@14693.4]
  wire  _T_1937; // @[package.scala 96:25:@14630.4 package.scala 96:25:@14631.4]
  wire  _T_2026; // @[package.scala 96:25:@14774.4 package.scala 96:25:@14775.4]
  wire [31:0] _T_2030; // @[Mux.scala 31:69:@14784.4]
  wire  _T_2023; // @[package.scala 96:25:@14766.4 package.scala 96:25:@14767.4]
  wire [31:0] _T_2031; // @[Mux.scala 31:69:@14785.4]
  wire  _T_2020; // @[package.scala 96:25:@14758.4 package.scala 96:25:@14759.4]
  wire [31:0] _T_2032; // @[Mux.scala 31:69:@14786.4]
  wire  _T_2017; // @[package.scala 96:25:@14750.4 package.scala 96:25:@14751.4]
  wire [31:0] _T_2033; // @[Mux.scala 31:69:@14787.4]
  wire  _T_2014; // @[package.scala 96:25:@14742.4 package.scala 96:25:@14743.4]
  wire [31:0] _T_2034; // @[Mux.scala 31:69:@14788.4]
  wire  _T_2011; // @[package.scala 96:25:@14734.4 package.scala 96:25:@14735.4]
  wire [31:0] _T_2035; // @[Mux.scala 31:69:@14789.4]
  wire  _T_2008; // @[package.scala 96:25:@14726.4 package.scala 96:25:@14727.4]
  wire  _T_2097; // @[package.scala 96:25:@14870.4 package.scala 96:25:@14871.4]
  wire [31:0] _T_2101; // @[Mux.scala 31:69:@14880.4]
  wire  _T_2094; // @[package.scala 96:25:@14862.4 package.scala 96:25:@14863.4]
  wire [31:0] _T_2102; // @[Mux.scala 31:69:@14881.4]
  wire  _T_2091; // @[package.scala 96:25:@14854.4 package.scala 96:25:@14855.4]
  wire [31:0] _T_2103; // @[Mux.scala 31:69:@14882.4]
  wire  _T_2088; // @[package.scala 96:25:@14846.4 package.scala 96:25:@14847.4]
  wire [31:0] _T_2104; // @[Mux.scala 31:69:@14883.4]
  wire  _T_2085; // @[package.scala 96:25:@14838.4 package.scala 96:25:@14839.4]
  wire [31:0] _T_2105; // @[Mux.scala 31:69:@14884.4]
  wire  _T_2082; // @[package.scala 96:25:@14830.4 package.scala 96:25:@14831.4]
  wire [31:0] _T_2106; // @[Mux.scala 31:69:@14885.4]
  wire  _T_2079; // @[package.scala 96:25:@14822.4 package.scala 96:25:@14823.4]
  wire  _T_2168; // @[package.scala 96:25:@14966.4 package.scala 96:25:@14967.4]
  wire [31:0] _T_2172; // @[Mux.scala 31:69:@14976.4]
  wire  _T_2165; // @[package.scala 96:25:@14958.4 package.scala 96:25:@14959.4]
  wire [31:0] _T_2173; // @[Mux.scala 31:69:@14977.4]
  wire  _T_2162; // @[package.scala 96:25:@14950.4 package.scala 96:25:@14951.4]
  wire [31:0] _T_2174; // @[Mux.scala 31:69:@14978.4]
  wire  _T_2159; // @[package.scala 96:25:@14942.4 package.scala 96:25:@14943.4]
  wire [31:0] _T_2175; // @[Mux.scala 31:69:@14979.4]
  wire  _T_2156; // @[package.scala 96:25:@14934.4 package.scala 96:25:@14935.4]
  wire [31:0] _T_2176; // @[Mux.scala 31:69:@14980.4]
  wire  _T_2153; // @[package.scala 96:25:@14926.4 package.scala 96:25:@14927.4]
  wire [31:0] _T_2177; // @[Mux.scala 31:69:@14981.4]
  wire  _T_2150; // @[package.scala 96:25:@14918.4 package.scala 96:25:@14919.4]
  wire  _T_2239; // @[package.scala 96:25:@15062.4 package.scala 96:25:@15063.4]
  wire [31:0] _T_2243; // @[Mux.scala 31:69:@15072.4]
  wire  _T_2236; // @[package.scala 96:25:@15054.4 package.scala 96:25:@15055.4]
  wire [31:0] _T_2244; // @[Mux.scala 31:69:@15073.4]
  wire  _T_2233; // @[package.scala 96:25:@15046.4 package.scala 96:25:@15047.4]
  wire [31:0] _T_2245; // @[Mux.scala 31:69:@15074.4]
  wire  _T_2230; // @[package.scala 96:25:@15038.4 package.scala 96:25:@15039.4]
  wire [31:0] _T_2246; // @[Mux.scala 31:69:@15075.4]
  wire  _T_2227; // @[package.scala 96:25:@15030.4 package.scala 96:25:@15031.4]
  wire [31:0] _T_2247; // @[Mux.scala 31:69:@15076.4]
  wire  _T_2224; // @[package.scala 96:25:@15022.4 package.scala 96:25:@15023.4]
  wire [31:0] _T_2248; // @[Mux.scala 31:69:@15077.4]
  wire  _T_2221; // @[package.scala 96:25:@15014.4 package.scala 96:25:@15015.4]
  wire  _T_2310; // @[package.scala 96:25:@15158.4 package.scala 96:25:@15159.4]
  wire [31:0] _T_2314; // @[Mux.scala 31:69:@15168.4]
  wire  _T_2307; // @[package.scala 96:25:@15150.4 package.scala 96:25:@15151.4]
  wire [31:0] _T_2315; // @[Mux.scala 31:69:@15169.4]
  wire  _T_2304; // @[package.scala 96:25:@15142.4 package.scala 96:25:@15143.4]
  wire [31:0] _T_2316; // @[Mux.scala 31:69:@15170.4]
  wire  _T_2301; // @[package.scala 96:25:@15134.4 package.scala 96:25:@15135.4]
  wire [31:0] _T_2317; // @[Mux.scala 31:69:@15171.4]
  wire  _T_2298; // @[package.scala 96:25:@15126.4 package.scala 96:25:@15127.4]
  wire [31:0] _T_2318; // @[Mux.scala 31:69:@15172.4]
  wire  _T_2295; // @[package.scala 96:25:@15118.4 package.scala 96:25:@15119.4]
  wire [31:0] _T_2319; // @[Mux.scala 31:69:@15173.4]
  wire  _T_2292; // @[package.scala 96:25:@15110.4 package.scala 96:25:@15111.4]
  wire  _T_2381; // @[package.scala 96:25:@15254.4 package.scala 96:25:@15255.4]
  wire [31:0] _T_2385; // @[Mux.scala 31:69:@15264.4]
  wire  _T_2378; // @[package.scala 96:25:@15246.4 package.scala 96:25:@15247.4]
  wire [31:0] _T_2386; // @[Mux.scala 31:69:@15265.4]
  wire  _T_2375; // @[package.scala 96:25:@15238.4 package.scala 96:25:@15239.4]
  wire [31:0] _T_2387; // @[Mux.scala 31:69:@15266.4]
  wire  _T_2372; // @[package.scala 96:25:@15230.4 package.scala 96:25:@15231.4]
  wire [31:0] _T_2388; // @[Mux.scala 31:69:@15267.4]
  wire  _T_2369; // @[package.scala 96:25:@15222.4 package.scala 96:25:@15223.4]
  wire [31:0] _T_2389; // @[Mux.scala 31:69:@15268.4]
  wire  _T_2366; // @[package.scala 96:25:@15214.4 package.scala 96:25:@15215.4]
  wire [31:0] _T_2390; // @[Mux.scala 31:69:@15269.4]
  wire  _T_2363; // @[package.scala 96:25:@15206.4 package.scala 96:25:@15207.4]
  wire  _T_2452; // @[package.scala 96:25:@15350.4 package.scala 96:25:@15351.4]
  wire [31:0] _T_2456; // @[Mux.scala 31:69:@15360.4]
  wire  _T_2449; // @[package.scala 96:25:@15342.4 package.scala 96:25:@15343.4]
  wire [31:0] _T_2457; // @[Mux.scala 31:69:@15361.4]
  wire  _T_2446; // @[package.scala 96:25:@15334.4 package.scala 96:25:@15335.4]
  wire [31:0] _T_2458; // @[Mux.scala 31:69:@15362.4]
  wire  _T_2443; // @[package.scala 96:25:@15326.4 package.scala 96:25:@15327.4]
  wire [31:0] _T_2459; // @[Mux.scala 31:69:@15363.4]
  wire  _T_2440; // @[package.scala 96:25:@15318.4 package.scala 96:25:@15319.4]
  wire [31:0] _T_2460; // @[Mux.scala 31:69:@15364.4]
  wire  _T_2437; // @[package.scala 96:25:@15310.4 package.scala 96:25:@15311.4]
  wire [31:0] _T_2461; // @[Mux.scala 31:69:@15365.4]
  wire  _T_2434; // @[package.scala 96:25:@15302.4 package.scala 96:25:@15303.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12776.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12792.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12808.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12824.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12840.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12856.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12872.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12888.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12904.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12920.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12936.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12952.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@12968.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@12984.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@13000.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@13016.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@13248.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@13310.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@13372.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13434.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13496.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13558.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13620.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13682.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13744.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13806.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13868.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@13930.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@13992.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@14054.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@14116.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@14178.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@14241.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@14249.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@14257.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@14265.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@14273.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@14281.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@14289.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@14297.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@14337.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@14345.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@14353.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14361.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14369.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14377.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14385.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14393.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14433.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14441.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14449.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14457.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14465.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14473.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14481.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14489.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14529.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14537.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14545.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14553.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14561.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14569.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14577.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14585.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14625.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14633.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14641.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14649.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14657.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14665.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14673.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14681.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14721.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14729.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14737.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14745.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14753.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14761.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14769.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14777.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14817.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14825.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14833.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14841.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14849.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14857.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14865.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14873.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14913.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14921.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14929.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14937.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14945.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14953.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14961.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14969.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@15009.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@15017.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@15025.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@15033.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@15041.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@15049.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@15057.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@15065.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@15105.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@15113.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@15121.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@15129.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@15137.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@15145.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@15153.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@15161.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@15201.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@15209.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@15217.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@15225.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@15233.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@15241.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@15249.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@15257.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@15297.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@15305.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@15313.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@15321.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@15329.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@15337.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15345.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15353.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13032.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@13033.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@13034.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@13035.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13037.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13044.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@13045.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@13046.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@13047.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13049.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@13057.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@13058.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@13059.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13061.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@13069.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@13070.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@13071.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13073.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13080.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@13082.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@13083.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13085.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13092.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@13094.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@13095.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13097.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@13106.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@13107.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13109.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@13118.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@13119.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13121.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13128.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@13130.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@13131.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13133.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13140.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@13142.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@13143.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13145.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@13154.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@13155.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13157.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@13166.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@13167.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13169.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13176.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@13178.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@13179.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13181.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13188.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@13190.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@13191.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13193.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@13202.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@13203.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13205.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@13214.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@13215.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13217.4]
  assign _T_620 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13224.4]
  assign _T_622 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13225.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@13226.4]
  assign _T_626 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13228.4]
  assign _T_628 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13229.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@13230.4]
  assign _T_632 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13232.4]
  assign _T_634 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13233.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@13234.4]
  assign _T_638 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13236.4]
  assign _T_640 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13237.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@13238.4]
  assign _T_644 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13240.4]
  assign _T_646 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13241.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@13242.4]
  assign _T_650 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13244.4]
  assign _T_652 = io_rPort_11_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13245.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@13246.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@13257.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@13258.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@13259.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@13260.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@13261.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@13262.4]
  assign _T_662 = {_T_655,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13264.4]
  assign _T_664 = {_T_656,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13266.4]
  assign _T_666 = {_T_657,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13268.4]
  assign _T_668 = {_T_658,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13270.4]
  assign _T_670 = {_T_659,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13272.4]
  assign _T_672 = {_T_660,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13274.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@13275.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@13276.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@13277.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@13278.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@13279.4]
  assign _T_682 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13286.4]
  assign _T_684 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13287.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_688 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13290.4]
  assign _T_690 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13291.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_694 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13294.4]
  assign _T_696 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13295.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@13296.4]
  assign _T_700 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13298.4]
  assign _T_702 = io_rPort_8_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13299.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@13300.4]
  assign _T_706 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13302.4]
  assign _T_708 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13303.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@13304.4]
  assign _T_712 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13306.4]
  assign _T_714 = io_rPort_10_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13307.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@13308.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@13319.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@13320.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@13321.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@13322.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@13323.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@13324.4]
  assign _T_724 = {_T_717,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13326.4]
  assign _T_726 = {_T_718,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13328.4]
  assign _T_728 = {_T_719,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13330.4]
  assign _T_730 = {_T_720,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13332.4]
  assign _T_732 = {_T_721,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13334.4]
  assign _T_734 = {_T_722,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13336.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@13337.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@13338.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@13339.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@13340.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@13341.4]
  assign _T_746 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13349.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@13350.4]
  assign _T_752 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13353.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@13354.4]
  assign _T_758 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13357.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@13358.4]
  assign _T_764 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13361.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@13362.4]
  assign _T_770 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13365.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@13366.4]
  assign _T_776 = io_rPort_11_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13369.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@13370.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@13381.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@13382.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@13383.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@13384.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@13385.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@13386.4]
  assign _T_786 = {_T_779,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13388.4]
  assign _T_788 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13390.4]
  assign _T_790 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13392.4]
  assign _T_792 = {_T_782,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13394.4]
  assign _T_794 = {_T_783,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13396.4]
  assign _T_796 = {_T_784,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13398.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@13399.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@13400.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@13401.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@13402.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@13403.4]
  assign _T_808 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13411.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@13412.4]
  assign _T_814 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13415.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@13416.4]
  assign _T_820 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13419.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@13420.4]
  assign _T_826 = io_rPort_8_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13423.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@13424.4]
  assign _T_832 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13427.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@13428.4]
  assign _T_838 = io_rPort_10_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13431.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@13432.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13443.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13444.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13445.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13446.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13447.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13448.4]
  assign _T_848 = {_T_841,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13450.4]
  assign _T_850 = {_T_842,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13452.4]
  assign _T_852 = {_T_843,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13454.4]
  assign _T_854 = {_T_844,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13456.4]
  assign _T_856 = {_T_845,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13458.4]
  assign _T_858 = {_T_846,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13460.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@13461.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@13462.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@13463.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@13464.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@13465.4]
  assign _T_868 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13472.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@13474.4]
  assign _T_874 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13476.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@13478.4]
  assign _T_880 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13480.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@13482.4]
  assign _T_886 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13484.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@13486.4]
  assign _T_892 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13488.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@13490.4]
  assign _T_898 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13492.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@13494.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13505.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13506.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13507.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13508.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13509.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13510.4]
  assign _T_910 = {_T_903,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13512.4]
  assign _T_912 = {_T_904,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13514.4]
  assign _T_914 = {_T_905,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13516.4]
  assign _T_916 = {_T_906,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13518.4]
  assign _T_918 = {_T_907,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13520.4]
  assign _T_920 = {_T_908,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13522.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@13523.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@13524.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@13525.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@13526.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@13527.4]
  assign _T_930 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13534.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@13536.4]
  assign _T_936 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13538.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@13540.4]
  assign _T_942 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13542.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@13544.4]
  assign _T_948 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13546.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@13548.4]
  assign _T_954 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13550.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@13552.4]
  assign _T_960 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13554.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@13556.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13567.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13568.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13569.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13570.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13571.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13572.4]
  assign _T_972 = {_T_965,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13574.4]
  assign _T_974 = {_T_966,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13576.4]
  assign _T_976 = {_T_967,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13578.4]
  assign _T_978 = {_T_968,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13580.4]
  assign _T_980 = {_T_969,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13582.4]
  assign _T_982 = {_T_970,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13584.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@13585.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@13586.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@13587.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@13588.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@13589.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@13598.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@13602.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@13606.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@13610.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@13614.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@13618.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13629.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13630.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13631.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13632.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13633.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13634.4]
  assign _T_1034 = {_T_1027,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13636.4]
  assign _T_1036 = {_T_1028,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13638.4]
  assign _T_1038 = {_T_1029,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13640.4]
  assign _T_1040 = {_T_1030,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13642.4]
  assign _T_1042 = {_T_1031,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13644.4]
  assign _T_1044 = {_T_1032,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13646.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@13647.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@13648.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@13649.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@13650.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@13651.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@13660.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@13664.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@13668.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@13672.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@13676.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@13680.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13691.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13692.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13693.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13694.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13695.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13696.4]
  assign _T_1096 = {_T_1089,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13698.4]
  assign _T_1098 = {_T_1090,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13700.4]
  assign _T_1100 = {_T_1091,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13702.4]
  assign _T_1102 = {_T_1092,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13704.4]
  assign _T_1104 = {_T_1093,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13706.4]
  assign _T_1106 = {_T_1094,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13708.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@13709.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@13710.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@13711.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@13712.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@13713.4]
  assign _T_1116 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13720.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@13722.4]
  assign _T_1122 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13724.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@13726.4]
  assign _T_1128 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13728.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@13730.4]
  assign _T_1134 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13732.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@13734.4]
  assign _T_1140 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13736.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@13738.4]
  assign _T_1146 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13740.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@13742.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13753.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13754.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13755.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13756.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13757.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13758.4]
  assign _T_1158 = {_T_1151,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13760.4]
  assign _T_1160 = {_T_1152,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13762.4]
  assign _T_1162 = {_T_1153,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13764.4]
  assign _T_1164 = {_T_1154,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13766.4]
  assign _T_1166 = {_T_1155,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13768.4]
  assign _T_1168 = {_T_1156,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13770.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@13771.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@13772.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@13773.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@13774.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@13775.4]
  assign _T_1178 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13782.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@13784.4]
  assign _T_1184 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13786.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@13788.4]
  assign _T_1190 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13790.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@13792.4]
  assign _T_1196 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13794.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@13796.4]
  assign _T_1202 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13798.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@13800.4]
  assign _T_1208 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13802.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@13804.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13815.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13816.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13817.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13818.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13819.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13820.4]
  assign _T_1220 = {_T_1213,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13822.4]
  assign _T_1222 = {_T_1214,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13824.4]
  assign _T_1224 = {_T_1215,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13826.4]
  assign _T_1226 = {_T_1216,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13828.4]
  assign _T_1228 = {_T_1217,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13830.4]
  assign _T_1230 = {_T_1218,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13832.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@13833.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@13834.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@13835.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@13836.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@13837.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@13846.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@13850.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@13854.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@13858.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@13862.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@13866.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13877.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13878.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13879.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13880.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13881.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13882.4]
  assign _T_1282 = {_T_1275,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13884.4]
  assign _T_1284 = {_T_1276,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13886.4]
  assign _T_1286 = {_T_1277,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13888.4]
  assign _T_1288 = {_T_1278,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13890.4]
  assign _T_1290 = {_T_1279,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13892.4]
  assign _T_1292 = {_T_1280,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13894.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@13895.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@13896.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@13897.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@13898.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@13899.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@13908.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@13912.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@13916.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@13920.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@13924.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@13928.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@13939.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@13940.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@13941.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@13942.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@13943.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@13944.4]
  assign _T_1344 = {_T_1337,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13946.4]
  assign _T_1346 = {_T_1338,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13948.4]
  assign _T_1348 = {_T_1339,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13950.4]
  assign _T_1350 = {_T_1340,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13952.4]
  assign _T_1352 = {_T_1341,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13954.4]
  assign _T_1354 = {_T_1342,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13956.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@13957.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@13958.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@13959.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@13960.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@13961.4]
  assign _T_1364 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13968.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@13970.4]
  assign _T_1370 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13972.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@13974.4]
  assign _T_1376 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13976.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@13978.4]
  assign _T_1382 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13980.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@13982.4]
  assign _T_1388 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13984.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@13986.4]
  assign _T_1394 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13988.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@13990.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@14001.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@14002.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@14003.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@14004.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@14005.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@14006.4]
  assign _T_1406 = {_T_1399,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14008.4]
  assign _T_1408 = {_T_1400,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14010.4]
  assign _T_1410 = {_T_1401,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14012.4]
  assign _T_1412 = {_T_1402,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14014.4]
  assign _T_1414 = {_T_1403,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14016.4]
  assign _T_1416 = {_T_1404,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@14018.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@14019.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@14020.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@14021.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@14022.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@14023.4]
  assign _T_1426 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14030.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@14032.4]
  assign _T_1432 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14034.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@14036.4]
  assign _T_1438 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14038.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@14040.4]
  assign _T_1444 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14042.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@14044.4]
  assign _T_1450 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14046.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@14048.4]
  assign _T_1456 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14050.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@14052.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@14063.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@14064.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@14065.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@14066.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@14067.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@14068.4]
  assign _T_1468 = {_T_1461,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14070.4]
  assign _T_1470 = {_T_1462,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14072.4]
  assign _T_1472 = {_T_1463,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14074.4]
  assign _T_1474 = {_T_1464,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14076.4]
  assign _T_1476 = {_T_1465,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14078.4]
  assign _T_1478 = {_T_1466,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@14080.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@14081.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@14082.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@14083.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@14084.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@14085.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@14094.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@14098.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@14102.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@14106.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@14110.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@14114.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@14125.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@14126.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@14127.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@14128.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@14129.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@14130.4]
  assign _T_1530 = {_T_1523,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14132.4]
  assign _T_1532 = {_T_1524,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14134.4]
  assign _T_1534 = {_T_1525,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14136.4]
  assign _T_1536 = {_T_1526,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14138.4]
  assign _T_1538 = {_T_1527,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14140.4]
  assign _T_1540 = {_T_1528,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@14142.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@14143.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@14144.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@14145.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@14146.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@14147.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@14156.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@14160.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@14164.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@14168.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@14172.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@14176.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@14187.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@14188.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@14189.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@14190.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@14191.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@14192.4]
  assign _T_1592 = {_T_1585,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14194.4]
  assign _T_1594 = {_T_1586,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14196.4]
  assign _T_1596 = {_T_1587,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14198.4]
  assign _T_1598 = {_T_1588,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14200.4]
  assign _T_1600 = {_T_1589,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14202.4]
  assign _T_1602 = {_T_1590,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@14204.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@14205.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@14206.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@14207.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@14208.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@14209.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14294.4 package.scala 96:25:@14295.4]
  assign _T_1675 = _T_1671 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14304.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14286.4 package.scala 96:25:@14287.4]
  assign _T_1676 = _T_1668 ? Mem1D_10_io_output : _T_1675; // @[Mux.scala 31:69:@14305.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14278.4 package.scala 96:25:@14279.4]
  assign _T_1677 = _T_1665 ? Mem1D_8_io_output : _T_1676; // @[Mux.scala 31:69:@14306.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14270.4 package.scala 96:25:@14271.4]
  assign _T_1678 = _T_1662 ? Mem1D_6_io_output : _T_1677; // @[Mux.scala 31:69:@14307.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14262.4 package.scala 96:25:@14263.4]
  assign _T_1679 = _T_1659 ? Mem1D_4_io_output : _T_1678; // @[Mux.scala 31:69:@14308.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14254.4 package.scala 96:25:@14255.4]
  assign _T_1680 = _T_1656 ? Mem1D_2_io_output : _T_1679; // @[Mux.scala 31:69:@14309.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@14246.4 package.scala 96:25:@14247.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14390.4 package.scala 96:25:@14391.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14400.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14382.4 package.scala 96:25:@14383.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@14401.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14374.4 package.scala 96:25:@14375.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@14402.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@14366.4 package.scala 96:25:@14367.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@14403.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14358.4 package.scala 96:25:@14359.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@14404.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14350.4 package.scala 96:25:@14351.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@14405.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14342.4 package.scala 96:25:@14343.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14486.4 package.scala 96:25:@14487.4]
  assign _T_1817 = _T_1813 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14496.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14478.4 package.scala 96:25:@14479.4]
  assign _T_1818 = _T_1810 ? Mem1D_11_io_output : _T_1817; // @[Mux.scala 31:69:@14497.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14470.4 package.scala 96:25:@14471.4]
  assign _T_1819 = _T_1807 ? Mem1D_9_io_output : _T_1818; // @[Mux.scala 31:69:@14498.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14462.4 package.scala 96:25:@14463.4]
  assign _T_1820 = _T_1804 ? Mem1D_7_io_output : _T_1819; // @[Mux.scala 31:69:@14499.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14454.4 package.scala 96:25:@14455.4]
  assign _T_1821 = _T_1801 ? Mem1D_5_io_output : _T_1820; // @[Mux.scala 31:69:@14500.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14446.4 package.scala 96:25:@14447.4]
  assign _T_1822 = _T_1798 ? Mem1D_3_io_output : _T_1821; // @[Mux.scala 31:69:@14501.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14438.4 package.scala 96:25:@14439.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14582.4 package.scala 96:25:@14583.4]
  assign _T_1888 = _T_1884 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14592.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14574.4 package.scala 96:25:@14575.4]
  assign _T_1889 = _T_1881 ? Mem1D_10_io_output : _T_1888; // @[Mux.scala 31:69:@14593.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14566.4 package.scala 96:25:@14567.4]
  assign _T_1890 = _T_1878 ? Mem1D_8_io_output : _T_1889; // @[Mux.scala 31:69:@14594.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14558.4 package.scala 96:25:@14559.4]
  assign _T_1891 = _T_1875 ? Mem1D_6_io_output : _T_1890; // @[Mux.scala 31:69:@14595.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14550.4 package.scala 96:25:@14551.4]
  assign _T_1892 = _T_1872 ? Mem1D_4_io_output : _T_1891; // @[Mux.scala 31:69:@14596.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14542.4 package.scala 96:25:@14543.4]
  assign _T_1893 = _T_1869 ? Mem1D_2_io_output : _T_1892; // @[Mux.scala 31:69:@14597.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14534.4 package.scala 96:25:@14535.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14678.4 package.scala 96:25:@14679.4]
  assign _T_1959 = _T_1955 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14688.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14670.4 package.scala 96:25:@14671.4]
  assign _T_1960 = _T_1952 ? Mem1D_10_io_output : _T_1959; // @[Mux.scala 31:69:@14689.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14662.4 package.scala 96:25:@14663.4]
  assign _T_1961 = _T_1949 ? Mem1D_8_io_output : _T_1960; // @[Mux.scala 31:69:@14690.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@14654.4 package.scala 96:25:@14655.4]
  assign _T_1962 = _T_1946 ? Mem1D_6_io_output : _T_1961; // @[Mux.scala 31:69:@14691.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14646.4 package.scala 96:25:@14647.4]
  assign _T_1963 = _T_1943 ? Mem1D_4_io_output : _T_1962; // @[Mux.scala 31:69:@14692.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14638.4 package.scala 96:25:@14639.4]
  assign _T_1964 = _T_1940 ? Mem1D_2_io_output : _T_1963; // @[Mux.scala 31:69:@14693.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14630.4 package.scala 96:25:@14631.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14774.4 package.scala 96:25:@14775.4]
  assign _T_2030 = _T_2026 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14784.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14766.4 package.scala 96:25:@14767.4]
  assign _T_2031 = _T_2023 ? Mem1D_11_io_output : _T_2030; // @[Mux.scala 31:69:@14785.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14758.4 package.scala 96:25:@14759.4]
  assign _T_2032 = _T_2020 ? Mem1D_9_io_output : _T_2031; // @[Mux.scala 31:69:@14786.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14750.4 package.scala 96:25:@14751.4]
  assign _T_2033 = _T_2017 ? Mem1D_7_io_output : _T_2032; // @[Mux.scala 31:69:@14787.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14742.4 package.scala 96:25:@14743.4]
  assign _T_2034 = _T_2014 ? Mem1D_5_io_output : _T_2033; // @[Mux.scala 31:69:@14788.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14734.4 package.scala 96:25:@14735.4]
  assign _T_2035 = _T_2011 ? Mem1D_3_io_output : _T_2034; // @[Mux.scala 31:69:@14789.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14726.4 package.scala 96:25:@14727.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14870.4 package.scala 96:25:@14871.4]
  assign _T_2101 = _T_2097 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14880.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14862.4 package.scala 96:25:@14863.4]
  assign _T_2102 = _T_2094 ? Mem1D_10_io_output : _T_2101; // @[Mux.scala 31:69:@14881.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14854.4 package.scala 96:25:@14855.4]
  assign _T_2103 = _T_2091 ? Mem1D_8_io_output : _T_2102; // @[Mux.scala 31:69:@14882.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14846.4 package.scala 96:25:@14847.4]
  assign _T_2104 = _T_2088 ? Mem1D_6_io_output : _T_2103; // @[Mux.scala 31:69:@14883.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14838.4 package.scala 96:25:@14839.4]
  assign _T_2105 = _T_2085 ? Mem1D_4_io_output : _T_2104; // @[Mux.scala 31:69:@14884.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14830.4 package.scala 96:25:@14831.4]
  assign _T_2106 = _T_2082 ? Mem1D_2_io_output : _T_2105; // @[Mux.scala 31:69:@14885.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14822.4 package.scala 96:25:@14823.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14966.4 package.scala 96:25:@14967.4]
  assign _T_2172 = _T_2168 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14976.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14958.4 package.scala 96:25:@14959.4]
  assign _T_2173 = _T_2165 ? Mem1D_10_io_output : _T_2172; // @[Mux.scala 31:69:@14977.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14950.4 package.scala 96:25:@14951.4]
  assign _T_2174 = _T_2162 ? Mem1D_8_io_output : _T_2173; // @[Mux.scala 31:69:@14978.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@14942.4 package.scala 96:25:@14943.4]
  assign _T_2175 = _T_2159 ? Mem1D_6_io_output : _T_2174; // @[Mux.scala 31:69:@14979.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14934.4 package.scala 96:25:@14935.4]
  assign _T_2176 = _T_2156 ? Mem1D_4_io_output : _T_2175; // @[Mux.scala 31:69:@14980.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14926.4 package.scala 96:25:@14927.4]
  assign _T_2177 = _T_2153 ? Mem1D_2_io_output : _T_2176; // @[Mux.scala 31:69:@14981.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14918.4 package.scala 96:25:@14919.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@15062.4 package.scala 96:25:@15063.4]
  assign _T_2243 = _T_2239 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15072.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@15054.4 package.scala 96:25:@15055.4]
  assign _T_2244 = _T_2236 ? Mem1D_11_io_output : _T_2243; // @[Mux.scala 31:69:@15073.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@15046.4 package.scala 96:25:@15047.4]
  assign _T_2245 = _T_2233 ? Mem1D_9_io_output : _T_2244; // @[Mux.scala 31:69:@15074.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@15038.4 package.scala 96:25:@15039.4]
  assign _T_2246 = _T_2230 ? Mem1D_7_io_output : _T_2245; // @[Mux.scala 31:69:@15075.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@15030.4 package.scala 96:25:@15031.4]
  assign _T_2247 = _T_2227 ? Mem1D_5_io_output : _T_2246; // @[Mux.scala 31:69:@15076.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@15022.4 package.scala 96:25:@15023.4]
  assign _T_2248 = _T_2224 ? Mem1D_3_io_output : _T_2247; // @[Mux.scala 31:69:@15077.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@15014.4 package.scala 96:25:@15015.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@15158.4 package.scala 96:25:@15159.4]
  assign _T_2314 = _T_2310 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15168.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@15150.4 package.scala 96:25:@15151.4]
  assign _T_2315 = _T_2307 ? Mem1D_11_io_output : _T_2314; // @[Mux.scala 31:69:@15169.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@15142.4 package.scala 96:25:@15143.4]
  assign _T_2316 = _T_2304 ? Mem1D_9_io_output : _T_2315; // @[Mux.scala 31:69:@15170.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@15134.4 package.scala 96:25:@15135.4]
  assign _T_2317 = _T_2301 ? Mem1D_7_io_output : _T_2316; // @[Mux.scala 31:69:@15171.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@15126.4 package.scala 96:25:@15127.4]
  assign _T_2318 = _T_2298 ? Mem1D_5_io_output : _T_2317; // @[Mux.scala 31:69:@15172.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@15118.4 package.scala 96:25:@15119.4]
  assign _T_2319 = _T_2295 ? Mem1D_3_io_output : _T_2318; // @[Mux.scala 31:69:@15173.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@15110.4 package.scala 96:25:@15111.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@15254.4 package.scala 96:25:@15255.4]
  assign _T_2385 = _T_2381 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15264.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@15246.4 package.scala 96:25:@15247.4]
  assign _T_2386 = _T_2378 ? Mem1D_11_io_output : _T_2385; // @[Mux.scala 31:69:@15265.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@15238.4 package.scala 96:25:@15239.4]
  assign _T_2387 = _T_2375 ? Mem1D_9_io_output : _T_2386; // @[Mux.scala 31:69:@15266.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@15230.4 package.scala 96:25:@15231.4]
  assign _T_2388 = _T_2372 ? Mem1D_7_io_output : _T_2387; // @[Mux.scala 31:69:@15267.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@15222.4 package.scala 96:25:@15223.4]
  assign _T_2389 = _T_2369 ? Mem1D_5_io_output : _T_2388; // @[Mux.scala 31:69:@15268.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@15214.4 package.scala 96:25:@15215.4]
  assign _T_2390 = _T_2366 ? Mem1D_3_io_output : _T_2389; // @[Mux.scala 31:69:@15269.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@15206.4 package.scala 96:25:@15207.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15350.4 package.scala 96:25:@15351.4]
  assign _T_2456 = _T_2452 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@15360.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15342.4 package.scala 96:25:@15343.4]
  assign _T_2457 = _T_2449 ? Mem1D_10_io_output : _T_2456; // @[Mux.scala 31:69:@15361.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@15334.4 package.scala 96:25:@15335.4]
  assign _T_2458 = _T_2446 ? Mem1D_8_io_output : _T_2457; // @[Mux.scala 31:69:@15362.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@15326.4 package.scala 96:25:@15327.4]
  assign _T_2459 = _T_2443 ? Mem1D_6_io_output : _T_2458; // @[Mux.scala 31:69:@15363.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@15318.4 package.scala 96:25:@15319.4]
  assign _T_2460 = _T_2440 ? Mem1D_4_io_output : _T_2459; // @[Mux.scala 31:69:@15364.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@15310.4 package.scala 96:25:@15311.4]
  assign _T_2461 = _T_2437 ? Mem1D_2_io_output : _T_2460; // @[Mux.scala 31:69:@15365.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@15302.4 package.scala 96:25:@15303.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_io_output : _T_2461; // @[MemPrimitives.scala 152:13:@15367.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_1_io_output : _T_2390; // @[MemPrimitives.scala 152:13:@15271.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_1_io_output : _T_2319; // @[MemPrimitives.scala 152:13:@15175.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_1_io_output : _T_2248; // @[MemPrimitives.scala 152:13:@15079.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_io_output : _T_2177; // @[MemPrimitives.scala 152:13:@14983.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_io_output : _T_2106; // @[MemPrimitives.scala 152:13:@14887.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_1_io_output : _T_2035; // @[MemPrimitives.scala 152:13:@14791.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_io_output : _T_1964; // @[MemPrimitives.scala 152:13:@14695.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_io_output : _T_1893; // @[MemPrimitives.scala 152:13:@14599.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_1_io_output : _T_1822; // @[MemPrimitives.scala 152:13:@14503.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 152:13:@14407.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_io_output : _T_1680; // @[MemPrimitives.scala 152:13:@14311.4]
  assign Mem1D_clock = clock; // @[:@12777.4]
  assign Mem1D_reset = reset; // @[:@12778.4]
  assign Mem1D_io_r_ofs_0 = _T_677[8:0]; // @[MemPrimitives.scala 131:28:@13283.4]
  assign Mem1D_io_r_backpressure = _T_677[9]; // @[MemPrimitives.scala 132:32:@13284.4]
  assign Mem1D_io_w_ofs_0 = _T_450[8:0]; // @[MemPrimitives.scala 94:28:@13041.4]
  assign Mem1D_io_w_data_0 = _T_450[40:9]; // @[MemPrimitives.scala 95:29:@13042.4]
  assign Mem1D_io_w_en_0 = _T_450[41]; // @[MemPrimitives.scala 96:27:@13043.4]
  assign Mem1D_1_clock = clock; // @[:@12793.4]
  assign Mem1D_1_reset = reset; // @[:@12794.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[8:0]; // @[MemPrimitives.scala 131:28:@13345.4]
  assign Mem1D_1_io_r_backpressure = _T_739[9]; // @[MemPrimitives.scala 132:32:@13346.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[8:0]; // @[MemPrimitives.scala 94:28:@13053.4]
  assign Mem1D_1_io_w_data_0 = _T_461[40:9]; // @[MemPrimitives.scala 95:29:@13054.4]
  assign Mem1D_1_io_w_en_0 = _T_461[41]; // @[MemPrimitives.scala 96:27:@13055.4]
  assign Mem1D_2_clock = clock; // @[:@12809.4]
  assign Mem1D_2_reset = reset; // @[:@12810.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[8:0]; // @[MemPrimitives.scala 131:28:@13407.4]
  assign Mem1D_2_io_r_backpressure = _T_801[9]; // @[MemPrimitives.scala 132:32:@13408.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[8:0]; // @[MemPrimitives.scala 94:28:@13065.4]
  assign Mem1D_2_io_w_data_0 = _T_472[40:9]; // @[MemPrimitives.scala 95:29:@13066.4]
  assign Mem1D_2_io_w_en_0 = _T_472[41]; // @[MemPrimitives.scala 96:27:@13067.4]
  assign Mem1D_3_clock = clock; // @[:@12825.4]
  assign Mem1D_3_reset = reset; // @[:@12826.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[8:0]; // @[MemPrimitives.scala 131:28:@13469.4]
  assign Mem1D_3_io_r_backpressure = _T_863[9]; // @[MemPrimitives.scala 132:32:@13470.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[8:0]; // @[MemPrimitives.scala 94:28:@13077.4]
  assign Mem1D_3_io_w_data_0 = _T_483[40:9]; // @[MemPrimitives.scala 95:29:@13078.4]
  assign Mem1D_3_io_w_en_0 = _T_483[41]; // @[MemPrimitives.scala 96:27:@13079.4]
  assign Mem1D_4_clock = clock; // @[:@12841.4]
  assign Mem1D_4_reset = reset; // @[:@12842.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[8:0]; // @[MemPrimitives.scala 131:28:@13531.4]
  assign Mem1D_4_io_r_backpressure = _T_925[9]; // @[MemPrimitives.scala 132:32:@13532.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[8:0]; // @[MemPrimitives.scala 94:28:@13089.4]
  assign Mem1D_4_io_w_data_0 = _T_494[40:9]; // @[MemPrimitives.scala 95:29:@13090.4]
  assign Mem1D_4_io_w_en_0 = _T_494[41]; // @[MemPrimitives.scala 96:27:@13091.4]
  assign Mem1D_5_clock = clock; // @[:@12857.4]
  assign Mem1D_5_reset = reset; // @[:@12858.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[8:0]; // @[MemPrimitives.scala 131:28:@13593.4]
  assign Mem1D_5_io_r_backpressure = _T_987[9]; // @[MemPrimitives.scala 132:32:@13594.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[8:0]; // @[MemPrimitives.scala 94:28:@13101.4]
  assign Mem1D_5_io_w_data_0 = _T_505[40:9]; // @[MemPrimitives.scala 95:29:@13102.4]
  assign Mem1D_5_io_w_en_0 = _T_505[41]; // @[MemPrimitives.scala 96:27:@13103.4]
  assign Mem1D_6_clock = clock; // @[:@12873.4]
  assign Mem1D_6_reset = reset; // @[:@12874.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[8:0]; // @[MemPrimitives.scala 131:28:@13655.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[9]; // @[MemPrimitives.scala 132:32:@13656.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[8:0]; // @[MemPrimitives.scala 94:28:@13113.4]
  assign Mem1D_6_io_w_data_0 = _T_516[40:9]; // @[MemPrimitives.scala 95:29:@13114.4]
  assign Mem1D_6_io_w_en_0 = _T_516[41]; // @[MemPrimitives.scala 96:27:@13115.4]
  assign Mem1D_7_clock = clock; // @[:@12889.4]
  assign Mem1D_7_reset = reset; // @[:@12890.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[8:0]; // @[MemPrimitives.scala 131:28:@13717.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[9]; // @[MemPrimitives.scala 132:32:@13718.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[8:0]; // @[MemPrimitives.scala 94:28:@13125.4]
  assign Mem1D_7_io_w_data_0 = _T_527[40:9]; // @[MemPrimitives.scala 95:29:@13126.4]
  assign Mem1D_7_io_w_en_0 = _T_527[41]; // @[MemPrimitives.scala 96:27:@13127.4]
  assign Mem1D_8_clock = clock; // @[:@12905.4]
  assign Mem1D_8_reset = reset; // @[:@12906.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[8:0]; // @[MemPrimitives.scala 131:28:@13779.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[9]; // @[MemPrimitives.scala 132:32:@13780.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[8:0]; // @[MemPrimitives.scala 94:28:@13137.4]
  assign Mem1D_8_io_w_data_0 = _T_538[40:9]; // @[MemPrimitives.scala 95:29:@13138.4]
  assign Mem1D_8_io_w_en_0 = _T_538[41]; // @[MemPrimitives.scala 96:27:@13139.4]
  assign Mem1D_9_clock = clock; // @[:@12921.4]
  assign Mem1D_9_reset = reset; // @[:@12922.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[8:0]; // @[MemPrimitives.scala 131:28:@13841.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[9]; // @[MemPrimitives.scala 132:32:@13842.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[8:0]; // @[MemPrimitives.scala 94:28:@13149.4]
  assign Mem1D_9_io_w_data_0 = _T_549[40:9]; // @[MemPrimitives.scala 95:29:@13150.4]
  assign Mem1D_9_io_w_en_0 = _T_549[41]; // @[MemPrimitives.scala 96:27:@13151.4]
  assign Mem1D_10_clock = clock; // @[:@12937.4]
  assign Mem1D_10_reset = reset; // @[:@12938.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[8:0]; // @[MemPrimitives.scala 131:28:@13903.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[9]; // @[MemPrimitives.scala 132:32:@13904.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[8:0]; // @[MemPrimitives.scala 94:28:@13161.4]
  assign Mem1D_10_io_w_data_0 = _T_560[40:9]; // @[MemPrimitives.scala 95:29:@13162.4]
  assign Mem1D_10_io_w_en_0 = _T_560[41]; // @[MemPrimitives.scala 96:27:@13163.4]
  assign Mem1D_11_clock = clock; // @[:@12953.4]
  assign Mem1D_11_reset = reset; // @[:@12954.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@13965.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@13966.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[8:0]; // @[MemPrimitives.scala 94:28:@13173.4]
  assign Mem1D_11_io_w_data_0 = _T_571[40:9]; // @[MemPrimitives.scala 95:29:@13174.4]
  assign Mem1D_11_io_w_en_0 = _T_571[41]; // @[MemPrimitives.scala 96:27:@13175.4]
  assign Mem1D_12_clock = clock; // @[:@12969.4]
  assign Mem1D_12_reset = reset; // @[:@12970.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[8:0]; // @[MemPrimitives.scala 131:28:@14027.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[9]; // @[MemPrimitives.scala 132:32:@14028.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[8:0]; // @[MemPrimitives.scala 94:28:@13185.4]
  assign Mem1D_12_io_w_data_0 = _T_582[40:9]; // @[MemPrimitives.scala 95:29:@13186.4]
  assign Mem1D_12_io_w_en_0 = _T_582[41]; // @[MemPrimitives.scala 96:27:@13187.4]
  assign Mem1D_13_clock = clock; // @[:@12985.4]
  assign Mem1D_13_reset = reset; // @[:@12986.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[8:0]; // @[MemPrimitives.scala 131:28:@14089.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[9]; // @[MemPrimitives.scala 132:32:@14090.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[8:0]; // @[MemPrimitives.scala 94:28:@13197.4]
  assign Mem1D_13_io_w_data_0 = _T_593[40:9]; // @[MemPrimitives.scala 95:29:@13198.4]
  assign Mem1D_13_io_w_en_0 = _T_593[41]; // @[MemPrimitives.scala 96:27:@13199.4]
  assign Mem1D_14_clock = clock; // @[:@13001.4]
  assign Mem1D_14_reset = reset; // @[:@13002.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[8:0]; // @[MemPrimitives.scala 131:28:@14151.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[9]; // @[MemPrimitives.scala 132:32:@14152.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[8:0]; // @[MemPrimitives.scala 94:28:@13209.4]
  assign Mem1D_14_io_w_data_0 = _T_604[40:9]; // @[MemPrimitives.scala 95:29:@13210.4]
  assign Mem1D_14_io_w_en_0 = _T_604[41]; // @[MemPrimitives.scala 96:27:@13211.4]
  assign Mem1D_15_clock = clock; // @[:@13017.4]
  assign Mem1D_15_reset = reset; // @[:@13018.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[8:0]; // @[MemPrimitives.scala 131:28:@14213.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[9]; // @[MemPrimitives.scala 132:32:@14214.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@13221.4]
  assign Mem1D_15_io_w_data_0 = _T_615[40:9]; // @[MemPrimitives.scala 95:29:@13222.4]
  assign Mem1D_15_io_w_en_0 = _T_615[41]; // @[MemPrimitives.scala 96:27:@13223.4]
  assign StickySelects_clock = clock; // @[:@13249.4]
  assign StickySelects_reset = reset; // @[:@13250.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_623; // @[MemPrimitives.scala 125:64:@13251.4]
  assign StickySelects_io_ins_1 = io_rPort_3_en_0 & _T_629; // @[MemPrimitives.scala 125:64:@13252.4]
  assign StickySelects_io_ins_2 = io_rPort_4_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@13253.4]
  assign StickySelects_io_ins_3 = io_rPort_6_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@13254.4]
  assign StickySelects_io_ins_4 = io_rPort_7_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@13255.4]
  assign StickySelects_io_ins_5 = io_rPort_11_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@13256.4]
  assign StickySelects_1_clock = clock; // @[:@13311.4]
  assign StickySelects_1_reset = reset; // @[:@13312.4]
  assign StickySelects_1_io_ins_0 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 125:64:@13313.4]
  assign StickySelects_1_io_ins_1 = io_rPort_2_en_0 & _T_691; // @[MemPrimitives.scala 125:64:@13314.4]
  assign StickySelects_1_io_ins_2 = io_rPort_5_en_0 & _T_697; // @[MemPrimitives.scala 125:64:@13315.4]
  assign StickySelects_1_io_ins_3 = io_rPort_8_en_0 & _T_703; // @[MemPrimitives.scala 125:64:@13316.4]
  assign StickySelects_1_io_ins_4 = io_rPort_9_en_0 & _T_709; // @[MemPrimitives.scala 125:64:@13317.4]
  assign StickySelects_1_io_ins_5 = io_rPort_10_en_0 & _T_715; // @[MemPrimitives.scala 125:64:@13318.4]
  assign StickySelects_2_clock = clock; // @[:@13373.4]
  assign StickySelects_2_reset = reset; // @[:@13374.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_747; // @[MemPrimitives.scala 125:64:@13375.4]
  assign StickySelects_2_io_ins_1 = io_rPort_3_en_0 & _T_753; // @[MemPrimitives.scala 125:64:@13376.4]
  assign StickySelects_2_io_ins_2 = io_rPort_4_en_0 & _T_759; // @[MemPrimitives.scala 125:64:@13377.4]
  assign StickySelects_2_io_ins_3 = io_rPort_6_en_0 & _T_765; // @[MemPrimitives.scala 125:64:@13378.4]
  assign StickySelects_2_io_ins_4 = io_rPort_7_en_0 & _T_771; // @[MemPrimitives.scala 125:64:@13379.4]
  assign StickySelects_2_io_ins_5 = io_rPort_11_en_0 & _T_777; // @[MemPrimitives.scala 125:64:@13380.4]
  assign StickySelects_3_clock = clock; // @[:@13435.4]
  assign StickySelects_3_reset = reset; // @[:@13436.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_809; // @[MemPrimitives.scala 125:64:@13437.4]
  assign StickySelects_3_io_ins_1 = io_rPort_2_en_0 & _T_815; // @[MemPrimitives.scala 125:64:@13438.4]
  assign StickySelects_3_io_ins_2 = io_rPort_5_en_0 & _T_821; // @[MemPrimitives.scala 125:64:@13439.4]
  assign StickySelects_3_io_ins_3 = io_rPort_8_en_0 & _T_827; // @[MemPrimitives.scala 125:64:@13440.4]
  assign StickySelects_3_io_ins_4 = io_rPort_9_en_0 & _T_833; // @[MemPrimitives.scala 125:64:@13441.4]
  assign StickySelects_3_io_ins_5 = io_rPort_10_en_0 & _T_839; // @[MemPrimitives.scala 125:64:@13442.4]
  assign StickySelects_4_clock = clock; // @[:@13497.4]
  assign StickySelects_4_reset = reset; // @[:@13498.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_871; // @[MemPrimitives.scala 125:64:@13499.4]
  assign StickySelects_4_io_ins_1 = io_rPort_3_en_0 & _T_877; // @[MemPrimitives.scala 125:64:@13500.4]
  assign StickySelects_4_io_ins_2 = io_rPort_4_en_0 & _T_883; // @[MemPrimitives.scala 125:64:@13501.4]
  assign StickySelects_4_io_ins_3 = io_rPort_6_en_0 & _T_889; // @[MemPrimitives.scala 125:64:@13502.4]
  assign StickySelects_4_io_ins_4 = io_rPort_7_en_0 & _T_895; // @[MemPrimitives.scala 125:64:@13503.4]
  assign StickySelects_4_io_ins_5 = io_rPort_11_en_0 & _T_901; // @[MemPrimitives.scala 125:64:@13504.4]
  assign StickySelects_5_clock = clock; // @[:@13559.4]
  assign StickySelects_5_reset = reset; // @[:@13560.4]
  assign StickySelects_5_io_ins_0 = io_rPort_1_en_0 & _T_933; // @[MemPrimitives.scala 125:64:@13561.4]
  assign StickySelects_5_io_ins_1 = io_rPort_2_en_0 & _T_939; // @[MemPrimitives.scala 125:64:@13562.4]
  assign StickySelects_5_io_ins_2 = io_rPort_5_en_0 & _T_945; // @[MemPrimitives.scala 125:64:@13563.4]
  assign StickySelects_5_io_ins_3 = io_rPort_8_en_0 & _T_951; // @[MemPrimitives.scala 125:64:@13564.4]
  assign StickySelects_5_io_ins_4 = io_rPort_9_en_0 & _T_957; // @[MemPrimitives.scala 125:64:@13565.4]
  assign StickySelects_5_io_ins_5 = io_rPort_10_en_0 & _T_963; // @[MemPrimitives.scala 125:64:@13566.4]
  assign StickySelects_6_clock = clock; // @[:@13621.4]
  assign StickySelects_6_reset = reset; // @[:@13622.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_995; // @[MemPrimitives.scala 125:64:@13623.4]
  assign StickySelects_6_io_ins_1 = io_rPort_3_en_0 & _T_1001; // @[MemPrimitives.scala 125:64:@13624.4]
  assign StickySelects_6_io_ins_2 = io_rPort_4_en_0 & _T_1007; // @[MemPrimitives.scala 125:64:@13625.4]
  assign StickySelects_6_io_ins_3 = io_rPort_6_en_0 & _T_1013; // @[MemPrimitives.scala 125:64:@13626.4]
  assign StickySelects_6_io_ins_4 = io_rPort_7_en_0 & _T_1019; // @[MemPrimitives.scala 125:64:@13627.4]
  assign StickySelects_6_io_ins_5 = io_rPort_11_en_0 & _T_1025; // @[MemPrimitives.scala 125:64:@13628.4]
  assign StickySelects_7_clock = clock; // @[:@13683.4]
  assign StickySelects_7_reset = reset; // @[:@13684.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1057; // @[MemPrimitives.scala 125:64:@13685.4]
  assign StickySelects_7_io_ins_1 = io_rPort_2_en_0 & _T_1063; // @[MemPrimitives.scala 125:64:@13686.4]
  assign StickySelects_7_io_ins_2 = io_rPort_5_en_0 & _T_1069; // @[MemPrimitives.scala 125:64:@13687.4]
  assign StickySelects_7_io_ins_3 = io_rPort_8_en_0 & _T_1075; // @[MemPrimitives.scala 125:64:@13688.4]
  assign StickySelects_7_io_ins_4 = io_rPort_9_en_0 & _T_1081; // @[MemPrimitives.scala 125:64:@13689.4]
  assign StickySelects_7_io_ins_5 = io_rPort_10_en_0 & _T_1087; // @[MemPrimitives.scala 125:64:@13690.4]
  assign StickySelects_8_clock = clock; // @[:@13745.4]
  assign StickySelects_8_reset = reset; // @[:@13746.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13747.4]
  assign StickySelects_8_io_ins_1 = io_rPort_3_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13748.4]
  assign StickySelects_8_io_ins_2 = io_rPort_4_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13749.4]
  assign StickySelects_8_io_ins_3 = io_rPort_6_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13750.4]
  assign StickySelects_8_io_ins_4 = io_rPort_7_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13751.4]
  assign StickySelects_8_io_ins_5 = io_rPort_11_en_0 & _T_1149; // @[MemPrimitives.scala 125:64:@13752.4]
  assign StickySelects_9_clock = clock; // @[:@13807.4]
  assign StickySelects_9_reset = reset; // @[:@13808.4]
  assign StickySelects_9_io_ins_0 = io_rPort_1_en_0 & _T_1181; // @[MemPrimitives.scala 125:64:@13809.4]
  assign StickySelects_9_io_ins_1 = io_rPort_2_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13810.4]
  assign StickySelects_9_io_ins_2 = io_rPort_5_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13811.4]
  assign StickySelects_9_io_ins_3 = io_rPort_8_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13812.4]
  assign StickySelects_9_io_ins_4 = io_rPort_9_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13813.4]
  assign StickySelects_9_io_ins_5 = io_rPort_10_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13814.4]
  assign StickySelects_10_clock = clock; // @[:@13869.4]
  assign StickySelects_10_reset = reset; // @[:@13870.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1243; // @[MemPrimitives.scala 125:64:@13871.4]
  assign StickySelects_10_io_ins_1 = io_rPort_3_en_0 & _T_1249; // @[MemPrimitives.scala 125:64:@13872.4]
  assign StickySelects_10_io_ins_2 = io_rPort_4_en_0 & _T_1255; // @[MemPrimitives.scala 125:64:@13873.4]
  assign StickySelects_10_io_ins_3 = io_rPort_6_en_0 & _T_1261; // @[MemPrimitives.scala 125:64:@13874.4]
  assign StickySelects_10_io_ins_4 = io_rPort_7_en_0 & _T_1267; // @[MemPrimitives.scala 125:64:@13875.4]
  assign StickySelects_10_io_ins_5 = io_rPort_11_en_0 & _T_1273; // @[MemPrimitives.scala 125:64:@13876.4]
  assign StickySelects_11_clock = clock; // @[:@13931.4]
  assign StickySelects_11_reset = reset; // @[:@13932.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@13933.4]
  assign StickySelects_11_io_ins_1 = io_rPort_2_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@13934.4]
  assign StickySelects_11_io_ins_2 = io_rPort_5_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@13935.4]
  assign StickySelects_11_io_ins_3 = io_rPort_8_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@13936.4]
  assign StickySelects_11_io_ins_4 = io_rPort_9_en_0 & _T_1329; // @[MemPrimitives.scala 125:64:@13937.4]
  assign StickySelects_11_io_ins_5 = io_rPort_10_en_0 & _T_1335; // @[MemPrimitives.scala 125:64:@13938.4]
  assign StickySelects_12_clock = clock; // @[:@13993.4]
  assign StickySelects_12_reset = reset; // @[:@13994.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@13995.4]
  assign StickySelects_12_io_ins_1 = io_rPort_3_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@13996.4]
  assign StickySelects_12_io_ins_2 = io_rPort_4_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@13997.4]
  assign StickySelects_12_io_ins_3 = io_rPort_6_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@13998.4]
  assign StickySelects_12_io_ins_4 = io_rPort_7_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@13999.4]
  assign StickySelects_12_io_ins_5 = io_rPort_11_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@14000.4]
  assign StickySelects_13_clock = clock; // @[:@14055.4]
  assign StickySelects_13_reset = reset; // @[:@14056.4]
  assign StickySelects_13_io_ins_0 = io_rPort_1_en_0 & _T_1429; // @[MemPrimitives.scala 125:64:@14057.4]
  assign StickySelects_13_io_ins_1 = io_rPort_2_en_0 & _T_1435; // @[MemPrimitives.scala 125:64:@14058.4]
  assign StickySelects_13_io_ins_2 = io_rPort_5_en_0 & _T_1441; // @[MemPrimitives.scala 125:64:@14059.4]
  assign StickySelects_13_io_ins_3 = io_rPort_8_en_0 & _T_1447; // @[MemPrimitives.scala 125:64:@14060.4]
  assign StickySelects_13_io_ins_4 = io_rPort_9_en_0 & _T_1453; // @[MemPrimitives.scala 125:64:@14061.4]
  assign StickySelects_13_io_ins_5 = io_rPort_10_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@14062.4]
  assign StickySelects_14_clock = clock; // @[:@14117.4]
  assign StickySelects_14_reset = reset; // @[:@14118.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_1491; // @[MemPrimitives.scala 125:64:@14119.4]
  assign StickySelects_14_io_ins_1 = io_rPort_3_en_0 & _T_1497; // @[MemPrimitives.scala 125:64:@14120.4]
  assign StickySelects_14_io_ins_2 = io_rPort_4_en_0 & _T_1503; // @[MemPrimitives.scala 125:64:@14121.4]
  assign StickySelects_14_io_ins_3 = io_rPort_6_en_0 & _T_1509; // @[MemPrimitives.scala 125:64:@14122.4]
  assign StickySelects_14_io_ins_4 = io_rPort_7_en_0 & _T_1515; // @[MemPrimitives.scala 125:64:@14123.4]
  assign StickySelects_14_io_ins_5 = io_rPort_11_en_0 & _T_1521; // @[MemPrimitives.scala 125:64:@14124.4]
  assign StickySelects_15_clock = clock; // @[:@14179.4]
  assign StickySelects_15_reset = reset; // @[:@14180.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_1553; // @[MemPrimitives.scala 125:64:@14181.4]
  assign StickySelects_15_io_ins_1 = io_rPort_2_en_0 & _T_1559; // @[MemPrimitives.scala 125:64:@14182.4]
  assign StickySelects_15_io_ins_2 = io_rPort_5_en_0 & _T_1565; // @[MemPrimitives.scala 125:64:@14183.4]
  assign StickySelects_15_io_ins_3 = io_rPort_8_en_0 & _T_1571; // @[MemPrimitives.scala 125:64:@14184.4]
  assign StickySelects_15_io_ins_4 = io_rPort_9_en_0 & _T_1577; // @[MemPrimitives.scala 125:64:@14185.4]
  assign StickySelects_15_io_ins_5 = io_rPort_10_en_0 & _T_1583; // @[MemPrimitives.scala 125:64:@14186.4]
  assign RetimeWrapper_clock = clock; // @[:@14242.4]
  assign RetimeWrapper_reset = reset; // @[:@14243.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14245.4]
  assign RetimeWrapper_io_in = _T_623 & io_rPort_0_en_0; // @[package.scala 94:16:@14244.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14250.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14251.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14253.4]
  assign RetimeWrapper_1_io_in = _T_747 & io_rPort_0_en_0; // @[package.scala 94:16:@14252.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14258.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14259.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14261.4]
  assign RetimeWrapper_2_io_in = _T_871 & io_rPort_0_en_0; // @[package.scala 94:16:@14260.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14266.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14267.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14269.4]
  assign RetimeWrapper_3_io_in = _T_995 & io_rPort_0_en_0; // @[package.scala 94:16:@14268.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14274.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14275.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14277.4]
  assign RetimeWrapper_4_io_in = _T_1119 & io_rPort_0_en_0; // @[package.scala 94:16:@14276.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14282.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14283.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14285.4]
  assign RetimeWrapper_5_io_in = _T_1243 & io_rPort_0_en_0; // @[package.scala 94:16:@14284.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14290.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14291.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14293.4]
  assign RetimeWrapper_6_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@14292.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14298.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14299.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14301.4]
  assign RetimeWrapper_7_io_in = _T_1491 & io_rPort_0_en_0; // @[package.scala 94:16:@14300.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14338.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14339.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14341.4]
  assign RetimeWrapper_8_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@14340.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14346.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14347.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14349.4]
  assign RetimeWrapper_9_io_in = _T_809 & io_rPort_1_en_0; // @[package.scala 94:16:@14348.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14354.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14355.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14357.4]
  assign RetimeWrapper_10_io_in = _T_933 & io_rPort_1_en_0; // @[package.scala 94:16:@14356.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14362.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14363.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14365.4]
  assign RetimeWrapper_11_io_in = _T_1057 & io_rPort_1_en_0; // @[package.scala 94:16:@14364.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14370.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14371.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14373.4]
  assign RetimeWrapper_12_io_in = _T_1181 & io_rPort_1_en_0; // @[package.scala 94:16:@14372.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14378.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14379.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14381.4]
  assign RetimeWrapper_13_io_in = _T_1305 & io_rPort_1_en_0; // @[package.scala 94:16:@14380.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14386.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14387.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14389.4]
  assign RetimeWrapper_14_io_in = _T_1429 & io_rPort_1_en_0; // @[package.scala 94:16:@14388.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14394.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14395.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14397.4]
  assign RetimeWrapper_15_io_in = _T_1553 & io_rPort_1_en_0; // @[package.scala 94:16:@14396.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14434.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14435.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14437.4]
  assign RetimeWrapper_16_io_in = _T_691 & io_rPort_2_en_0; // @[package.scala 94:16:@14436.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14442.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14443.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14445.4]
  assign RetimeWrapper_17_io_in = _T_815 & io_rPort_2_en_0; // @[package.scala 94:16:@14444.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14450.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14451.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14453.4]
  assign RetimeWrapper_18_io_in = _T_939 & io_rPort_2_en_0; // @[package.scala 94:16:@14452.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14458.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14459.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14461.4]
  assign RetimeWrapper_19_io_in = _T_1063 & io_rPort_2_en_0; // @[package.scala 94:16:@14460.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14466.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14467.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14469.4]
  assign RetimeWrapper_20_io_in = _T_1187 & io_rPort_2_en_0; // @[package.scala 94:16:@14468.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14474.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14475.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14477.4]
  assign RetimeWrapper_21_io_in = _T_1311 & io_rPort_2_en_0; // @[package.scala 94:16:@14476.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14482.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14483.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14485.4]
  assign RetimeWrapper_22_io_in = _T_1435 & io_rPort_2_en_0; // @[package.scala 94:16:@14484.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14490.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14491.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14493.4]
  assign RetimeWrapper_23_io_in = _T_1559 & io_rPort_2_en_0; // @[package.scala 94:16:@14492.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14530.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14531.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14533.4]
  assign RetimeWrapper_24_io_in = _T_629 & io_rPort_3_en_0; // @[package.scala 94:16:@14532.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14538.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14539.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14541.4]
  assign RetimeWrapper_25_io_in = _T_753 & io_rPort_3_en_0; // @[package.scala 94:16:@14540.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14546.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14547.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14549.4]
  assign RetimeWrapper_26_io_in = _T_877 & io_rPort_3_en_0; // @[package.scala 94:16:@14548.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14554.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14555.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14557.4]
  assign RetimeWrapper_27_io_in = _T_1001 & io_rPort_3_en_0; // @[package.scala 94:16:@14556.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14562.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14563.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14565.4]
  assign RetimeWrapper_28_io_in = _T_1125 & io_rPort_3_en_0; // @[package.scala 94:16:@14564.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14570.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14571.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14573.4]
  assign RetimeWrapper_29_io_in = _T_1249 & io_rPort_3_en_0; // @[package.scala 94:16:@14572.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14578.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14579.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14581.4]
  assign RetimeWrapper_30_io_in = _T_1373 & io_rPort_3_en_0; // @[package.scala 94:16:@14580.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14586.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14587.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14589.4]
  assign RetimeWrapper_31_io_in = _T_1497 & io_rPort_3_en_0; // @[package.scala 94:16:@14588.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14626.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14627.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14629.4]
  assign RetimeWrapper_32_io_in = _T_635 & io_rPort_4_en_0; // @[package.scala 94:16:@14628.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14634.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14635.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14637.4]
  assign RetimeWrapper_33_io_in = _T_759 & io_rPort_4_en_0; // @[package.scala 94:16:@14636.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14642.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14643.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14645.4]
  assign RetimeWrapper_34_io_in = _T_883 & io_rPort_4_en_0; // @[package.scala 94:16:@14644.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14650.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14651.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14653.4]
  assign RetimeWrapper_35_io_in = _T_1007 & io_rPort_4_en_0; // @[package.scala 94:16:@14652.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14658.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14659.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14661.4]
  assign RetimeWrapper_36_io_in = _T_1131 & io_rPort_4_en_0; // @[package.scala 94:16:@14660.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14666.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14667.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14669.4]
  assign RetimeWrapper_37_io_in = _T_1255 & io_rPort_4_en_0; // @[package.scala 94:16:@14668.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14674.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14675.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14677.4]
  assign RetimeWrapper_38_io_in = _T_1379 & io_rPort_4_en_0; // @[package.scala 94:16:@14676.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14682.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14683.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14685.4]
  assign RetimeWrapper_39_io_in = _T_1503 & io_rPort_4_en_0; // @[package.scala 94:16:@14684.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14722.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14723.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14725.4]
  assign RetimeWrapper_40_io_in = _T_697 & io_rPort_5_en_0; // @[package.scala 94:16:@14724.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14730.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14731.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14733.4]
  assign RetimeWrapper_41_io_in = _T_821 & io_rPort_5_en_0; // @[package.scala 94:16:@14732.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14738.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14739.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14741.4]
  assign RetimeWrapper_42_io_in = _T_945 & io_rPort_5_en_0; // @[package.scala 94:16:@14740.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14746.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14747.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14749.4]
  assign RetimeWrapper_43_io_in = _T_1069 & io_rPort_5_en_0; // @[package.scala 94:16:@14748.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14754.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14755.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14757.4]
  assign RetimeWrapper_44_io_in = _T_1193 & io_rPort_5_en_0; // @[package.scala 94:16:@14756.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14762.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14763.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14765.4]
  assign RetimeWrapper_45_io_in = _T_1317 & io_rPort_5_en_0; // @[package.scala 94:16:@14764.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14770.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14771.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14773.4]
  assign RetimeWrapper_46_io_in = _T_1441 & io_rPort_5_en_0; // @[package.scala 94:16:@14772.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14778.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14779.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14781.4]
  assign RetimeWrapper_47_io_in = _T_1565 & io_rPort_5_en_0; // @[package.scala 94:16:@14780.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14818.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14819.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14821.4]
  assign RetimeWrapper_48_io_in = _T_641 & io_rPort_6_en_0; // @[package.scala 94:16:@14820.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14826.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14827.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14829.4]
  assign RetimeWrapper_49_io_in = _T_765 & io_rPort_6_en_0; // @[package.scala 94:16:@14828.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14834.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14835.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14837.4]
  assign RetimeWrapper_50_io_in = _T_889 & io_rPort_6_en_0; // @[package.scala 94:16:@14836.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14842.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14843.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14845.4]
  assign RetimeWrapper_51_io_in = _T_1013 & io_rPort_6_en_0; // @[package.scala 94:16:@14844.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14850.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14851.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14853.4]
  assign RetimeWrapper_52_io_in = _T_1137 & io_rPort_6_en_0; // @[package.scala 94:16:@14852.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14858.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14859.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14861.4]
  assign RetimeWrapper_53_io_in = _T_1261 & io_rPort_6_en_0; // @[package.scala 94:16:@14860.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14866.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14867.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14869.4]
  assign RetimeWrapper_54_io_in = _T_1385 & io_rPort_6_en_0; // @[package.scala 94:16:@14868.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14874.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14875.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14877.4]
  assign RetimeWrapper_55_io_in = _T_1509 & io_rPort_6_en_0; // @[package.scala 94:16:@14876.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14914.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14915.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14917.4]
  assign RetimeWrapper_56_io_in = _T_647 & io_rPort_7_en_0; // @[package.scala 94:16:@14916.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14922.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14923.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14925.4]
  assign RetimeWrapper_57_io_in = _T_771 & io_rPort_7_en_0; // @[package.scala 94:16:@14924.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14930.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14931.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14933.4]
  assign RetimeWrapper_58_io_in = _T_895 & io_rPort_7_en_0; // @[package.scala 94:16:@14932.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14938.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14939.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14941.4]
  assign RetimeWrapper_59_io_in = _T_1019 & io_rPort_7_en_0; // @[package.scala 94:16:@14940.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14946.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14947.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14949.4]
  assign RetimeWrapper_60_io_in = _T_1143 & io_rPort_7_en_0; // @[package.scala 94:16:@14948.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14954.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14955.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14957.4]
  assign RetimeWrapper_61_io_in = _T_1267 & io_rPort_7_en_0; // @[package.scala 94:16:@14956.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14962.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14963.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14965.4]
  assign RetimeWrapper_62_io_in = _T_1391 & io_rPort_7_en_0; // @[package.scala 94:16:@14964.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14970.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14971.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14973.4]
  assign RetimeWrapper_63_io_in = _T_1515 & io_rPort_7_en_0; // @[package.scala 94:16:@14972.4]
  assign RetimeWrapper_64_clock = clock; // @[:@15010.4]
  assign RetimeWrapper_64_reset = reset; // @[:@15011.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15013.4]
  assign RetimeWrapper_64_io_in = _T_703 & io_rPort_8_en_0; // @[package.scala 94:16:@15012.4]
  assign RetimeWrapper_65_clock = clock; // @[:@15018.4]
  assign RetimeWrapper_65_reset = reset; // @[:@15019.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15021.4]
  assign RetimeWrapper_65_io_in = _T_827 & io_rPort_8_en_0; // @[package.scala 94:16:@15020.4]
  assign RetimeWrapper_66_clock = clock; // @[:@15026.4]
  assign RetimeWrapper_66_reset = reset; // @[:@15027.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15029.4]
  assign RetimeWrapper_66_io_in = _T_951 & io_rPort_8_en_0; // @[package.scala 94:16:@15028.4]
  assign RetimeWrapper_67_clock = clock; // @[:@15034.4]
  assign RetimeWrapper_67_reset = reset; // @[:@15035.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15037.4]
  assign RetimeWrapper_67_io_in = _T_1075 & io_rPort_8_en_0; // @[package.scala 94:16:@15036.4]
  assign RetimeWrapper_68_clock = clock; // @[:@15042.4]
  assign RetimeWrapper_68_reset = reset; // @[:@15043.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15045.4]
  assign RetimeWrapper_68_io_in = _T_1199 & io_rPort_8_en_0; // @[package.scala 94:16:@15044.4]
  assign RetimeWrapper_69_clock = clock; // @[:@15050.4]
  assign RetimeWrapper_69_reset = reset; // @[:@15051.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15053.4]
  assign RetimeWrapper_69_io_in = _T_1323 & io_rPort_8_en_0; // @[package.scala 94:16:@15052.4]
  assign RetimeWrapper_70_clock = clock; // @[:@15058.4]
  assign RetimeWrapper_70_reset = reset; // @[:@15059.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15061.4]
  assign RetimeWrapper_70_io_in = _T_1447 & io_rPort_8_en_0; // @[package.scala 94:16:@15060.4]
  assign RetimeWrapper_71_clock = clock; // @[:@15066.4]
  assign RetimeWrapper_71_reset = reset; // @[:@15067.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15069.4]
  assign RetimeWrapper_71_io_in = _T_1571 & io_rPort_8_en_0; // @[package.scala 94:16:@15068.4]
  assign RetimeWrapper_72_clock = clock; // @[:@15106.4]
  assign RetimeWrapper_72_reset = reset; // @[:@15107.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15109.4]
  assign RetimeWrapper_72_io_in = _T_709 & io_rPort_9_en_0; // @[package.scala 94:16:@15108.4]
  assign RetimeWrapper_73_clock = clock; // @[:@15114.4]
  assign RetimeWrapper_73_reset = reset; // @[:@15115.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15117.4]
  assign RetimeWrapper_73_io_in = _T_833 & io_rPort_9_en_0; // @[package.scala 94:16:@15116.4]
  assign RetimeWrapper_74_clock = clock; // @[:@15122.4]
  assign RetimeWrapper_74_reset = reset; // @[:@15123.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15125.4]
  assign RetimeWrapper_74_io_in = _T_957 & io_rPort_9_en_0; // @[package.scala 94:16:@15124.4]
  assign RetimeWrapper_75_clock = clock; // @[:@15130.4]
  assign RetimeWrapper_75_reset = reset; // @[:@15131.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15133.4]
  assign RetimeWrapper_75_io_in = _T_1081 & io_rPort_9_en_0; // @[package.scala 94:16:@15132.4]
  assign RetimeWrapper_76_clock = clock; // @[:@15138.4]
  assign RetimeWrapper_76_reset = reset; // @[:@15139.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15141.4]
  assign RetimeWrapper_76_io_in = _T_1205 & io_rPort_9_en_0; // @[package.scala 94:16:@15140.4]
  assign RetimeWrapper_77_clock = clock; // @[:@15146.4]
  assign RetimeWrapper_77_reset = reset; // @[:@15147.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15149.4]
  assign RetimeWrapper_77_io_in = _T_1329 & io_rPort_9_en_0; // @[package.scala 94:16:@15148.4]
  assign RetimeWrapper_78_clock = clock; // @[:@15154.4]
  assign RetimeWrapper_78_reset = reset; // @[:@15155.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15157.4]
  assign RetimeWrapper_78_io_in = _T_1453 & io_rPort_9_en_0; // @[package.scala 94:16:@15156.4]
  assign RetimeWrapper_79_clock = clock; // @[:@15162.4]
  assign RetimeWrapper_79_reset = reset; // @[:@15163.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15165.4]
  assign RetimeWrapper_79_io_in = _T_1577 & io_rPort_9_en_0; // @[package.scala 94:16:@15164.4]
  assign RetimeWrapper_80_clock = clock; // @[:@15202.4]
  assign RetimeWrapper_80_reset = reset; // @[:@15203.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15205.4]
  assign RetimeWrapper_80_io_in = _T_715 & io_rPort_10_en_0; // @[package.scala 94:16:@15204.4]
  assign RetimeWrapper_81_clock = clock; // @[:@15210.4]
  assign RetimeWrapper_81_reset = reset; // @[:@15211.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15213.4]
  assign RetimeWrapper_81_io_in = _T_839 & io_rPort_10_en_0; // @[package.scala 94:16:@15212.4]
  assign RetimeWrapper_82_clock = clock; // @[:@15218.4]
  assign RetimeWrapper_82_reset = reset; // @[:@15219.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15221.4]
  assign RetimeWrapper_82_io_in = _T_963 & io_rPort_10_en_0; // @[package.scala 94:16:@15220.4]
  assign RetimeWrapper_83_clock = clock; // @[:@15226.4]
  assign RetimeWrapper_83_reset = reset; // @[:@15227.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15229.4]
  assign RetimeWrapper_83_io_in = _T_1087 & io_rPort_10_en_0; // @[package.scala 94:16:@15228.4]
  assign RetimeWrapper_84_clock = clock; // @[:@15234.4]
  assign RetimeWrapper_84_reset = reset; // @[:@15235.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15237.4]
  assign RetimeWrapper_84_io_in = _T_1211 & io_rPort_10_en_0; // @[package.scala 94:16:@15236.4]
  assign RetimeWrapper_85_clock = clock; // @[:@15242.4]
  assign RetimeWrapper_85_reset = reset; // @[:@15243.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15245.4]
  assign RetimeWrapper_85_io_in = _T_1335 & io_rPort_10_en_0; // @[package.scala 94:16:@15244.4]
  assign RetimeWrapper_86_clock = clock; // @[:@15250.4]
  assign RetimeWrapper_86_reset = reset; // @[:@15251.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15253.4]
  assign RetimeWrapper_86_io_in = _T_1459 & io_rPort_10_en_0; // @[package.scala 94:16:@15252.4]
  assign RetimeWrapper_87_clock = clock; // @[:@15258.4]
  assign RetimeWrapper_87_reset = reset; // @[:@15259.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15261.4]
  assign RetimeWrapper_87_io_in = _T_1583 & io_rPort_10_en_0; // @[package.scala 94:16:@15260.4]
  assign RetimeWrapper_88_clock = clock; // @[:@15298.4]
  assign RetimeWrapper_88_reset = reset; // @[:@15299.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15301.4]
  assign RetimeWrapper_88_io_in = _T_653 & io_rPort_11_en_0; // @[package.scala 94:16:@15300.4]
  assign RetimeWrapper_89_clock = clock; // @[:@15306.4]
  assign RetimeWrapper_89_reset = reset; // @[:@15307.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15309.4]
  assign RetimeWrapper_89_io_in = _T_777 & io_rPort_11_en_0; // @[package.scala 94:16:@15308.4]
  assign RetimeWrapper_90_clock = clock; // @[:@15314.4]
  assign RetimeWrapper_90_reset = reset; // @[:@15315.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15317.4]
  assign RetimeWrapper_90_io_in = _T_901 & io_rPort_11_en_0; // @[package.scala 94:16:@15316.4]
  assign RetimeWrapper_91_clock = clock; // @[:@15322.4]
  assign RetimeWrapper_91_reset = reset; // @[:@15323.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15325.4]
  assign RetimeWrapper_91_io_in = _T_1025 & io_rPort_11_en_0; // @[package.scala 94:16:@15324.4]
  assign RetimeWrapper_92_clock = clock; // @[:@15330.4]
  assign RetimeWrapper_92_reset = reset; // @[:@15331.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15333.4]
  assign RetimeWrapper_92_io_in = _T_1149 & io_rPort_11_en_0; // @[package.scala 94:16:@15332.4]
  assign RetimeWrapper_93_clock = clock; // @[:@15338.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15339.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15341.4]
  assign RetimeWrapper_93_io_in = _T_1273 & io_rPort_11_en_0; // @[package.scala 94:16:@15340.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15346.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15347.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15349.4]
  assign RetimeWrapper_94_io_in = _T_1397 & io_rPort_11_en_0; // @[package.scala 94:16:@15348.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15354.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15355.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15357.4]
  assign RetimeWrapper_95_io_in = _T_1521 & io_rPort_11_en_0; // @[package.scala 94:16:@15356.4]
endmodule
module RetimeWrapper_168( // @[:@15772.2]
  input         clock, // @[:@15773.4]
  input         reset, // @[:@15774.4]
  input         io_flow, // @[:@15775.4]
  input  [31:0] io_in, // @[:@15775.4]
  output [31:0] io_out // @[:@15775.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15777.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15790.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15789.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15788.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15787.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15786.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15784.4]
endmodule
module RetimeWrapper_169( // @[:@15804.2]
  input   clock, // @[:@15805.4]
  input   reset, // @[:@15806.4]
  input   io_flow, // @[:@15807.4]
  input   io_in, // @[:@15807.4]
  output  io_out // @[:@15807.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15809.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15822.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15821.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15820.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15819.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15818.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15816.4]
endmodule
module RetimeWrapper_170( // @[:@15836.2]
  input         clock, // @[:@15837.4]
  input         reset, // @[:@15838.4]
  input         io_flow, // @[:@15839.4]
  input  [31:0] io_in, // @[:@15839.4]
  output [31:0] io_out // @[:@15839.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@15841.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15854.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15853.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15852.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15851.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15850.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15848.4]
endmodule
module RetimeWrapper_181( // @[:@16482.2]
  input         clock, // @[:@16483.4]
  input         reset, // @[:@16484.4]
  input         io_flow, // @[:@16485.4]
  input  [31:0] io_in, // @[:@16485.4]
  output [31:0] io_out // @[:@16485.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@16487.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16500.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16499.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16498.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16497.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16496.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16494.4]
endmodule
module RetimeWrapper_184( // @[:@16578.2]
  input         clock, // @[:@16579.4]
  input         reset, // @[:@16580.4]
  input         io_flow, // @[:@16581.4]
  input  [31:0] io_in, // @[:@16581.4]
  output [31:0] io_out // @[:@16581.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@16583.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16596.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16595.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16594.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16593.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16592.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16590.4]
endmodule
module RetimeWrapper_185( // @[:@16610.2]
  input         clock, // @[:@16611.4]
  input         reset, // @[:@16612.4]
  input         io_flow, // @[:@16613.4]
  input  [31:0] io_in, // @[:@16613.4]
  output [31:0] io_out // @[:@16613.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16615.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16615.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16615.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16615.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16615.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16615.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@16615.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16628.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16627.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16626.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16625.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16624.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16622.4]
endmodule
module RetimeWrapper_186( // @[:@16642.2]
  input   clock, // @[:@16643.4]
  input   reset, // @[:@16644.4]
  input   io_flow, // @[:@16645.4]
  input   io_in, // @[:@16645.4]
  output  io_out // @[:@16645.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@16647.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16660.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16659.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@16658.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16657.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16656.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16654.4]
endmodule
module RetimeWrapper_189( // @[:@16738.2]
  input         clock, // @[:@16739.4]
  input         reset, // @[:@16740.4]
  input         io_flow, // @[:@16741.4]
  input  [31:0] io_in, // @[:@16741.4]
  output [31:0] io_out // @[:@16741.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@16743.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16756.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16755.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16754.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16753.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16752.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16750.4]
endmodule
module Multiplier( // @[:@20852.2]
  input         clock, // @[:@20853.4]
  input         io_flow, // @[:@20855.4]
  input  [31:0] io_a, // @[:@20855.4]
  input  [31:0] io_b, // @[:@20855.4]
  output [31:0] io_out // @[:@20855.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@20857.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@20867.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@20865.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@20864.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@20866.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@20863.4]
endmodule
module x377( // @[:@20887.2]
  input         clock, // @[:@20888.4]
  input  [31:0] io_a, // @[:@20890.4]
  input  [31:0] io_b, // @[:@20890.4]
  input         io_flow, // @[:@20890.4]
  output [31:0] io_result // @[:@20890.4]
);
  wire  x377_clock; // @[BigIPZynq.scala 63:21:@20897.4]
  wire  x377_io_flow; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] x377_io_a; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] x377_io_b; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] x377_io_out; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@20906.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@20906.4]
  Multiplier x377 ( // @[BigIPZynq.scala 63:21:@20897.4]
    .clock(x377_clock),
    .io_flow(x377_io_flow),
    .io_a(x377_io_a),
    .io_b(x377_io_b),
    .io_out(x377_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@20906.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@20914.4]
  assign x377_clock = clock; // @[:@20898.4]
  assign x377_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@20902.4]
  assign x377_io_a = io_a; // @[BigIPZynq.scala 64:14:@20900.4]
  assign x377_io_b = io_b; // @[BigIPZynq.scala 65:14:@20901.4]
  assign fix2fixBox_io_a = x377_io_out; // @[Math.scala 254:23:@20909.4]
endmodule
module fix2fixBox_93( // @[:@21508.2]
  input  [31:0] io_a, // @[:@21511.4]
  output [32:0] io_b // @[:@21511.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@21525.4]
endmodule
module __56( // @[:@21527.2]
  input  [31:0] io_b, // @[:@21530.4]
  output [32:0] io_result // @[:@21530.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@21535.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@21535.4]
  fix2fixBox_93 fix2fixBox ( // @[BigIPZynq.scala 219:30:@21535.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@21543.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@21538.4]
endmodule
module x386_x13( // @[:@21639.2]
  input         clock, // @[:@21640.4]
  input         reset, // @[:@21641.4]
  input  [31:0] io_a, // @[:@21642.4]
  input  [31:0] io_b, // @[:@21642.4]
  input         io_flow, // @[:@21642.4]
  output [31:0] io_result // @[:@21642.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@21650.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@21650.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@21657.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@21657.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@21667.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@21667.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@21667.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@21667.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@21667.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@21655.4 Math.scala 724:14:@21656.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@21662.4 Math.scala 724:14:@21663.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@21664.4]
  __56 _ ( // @[Math.scala 720:24:@21650.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __56 __1 ( // @[Math.scala 720:24:@21657.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@21667.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@21655.4 Math.scala 724:14:@21656.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@21662.4 Math.scala 724:14:@21663.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@21664.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@21675.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@21653.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@21660.4]
  assign fix2fixBox_clock = clock; // @[:@21668.4]
  assign fix2fixBox_reset = reset; // @[:@21669.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@21670.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@21673.4]
endmodule
module fix2fixBox_117( // @[:@22892.2]
  input  [31:0] io_a, // @[:@22895.4]
  output [31:0] io_b // @[:@22895.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@22905.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@22905.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@22908.4]
endmodule
module x394( // @[:@22910.2]
  input  [31:0] io_b, // @[:@22913.4]
  output [31:0] io_result // @[:@22913.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@22918.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@22918.4]
  fix2fixBox_117 fix2fixBox ( // @[BigIPZynq.scala 219:30:@22918.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@22926.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@22921.4]
endmodule
module Multiplier_9( // @[:@22938.2]
  input         clock, // @[:@22939.4]
  input         io_flow, // @[:@22941.4]
  input  [38:0] io_a, // @[:@22941.4]
  input  [38:0] io_b, // @[:@22941.4]
  output [38:0] io_out // @[:@22941.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@22943.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@22953.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@22951.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@22950.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@22952.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@22949.4]
endmodule
module fix2fixBox_118( // @[:@22955.2]
  input  [38:0] io_a, // @[:@22958.4]
  output [31:0] io_b // @[:@22958.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@22966.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@22969.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@22966.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@22969.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@22972.4]
endmodule
module x395_mul( // @[:@22974.2]
  input         clock, // @[:@22975.4]
  input  [31:0] io_a, // @[:@22977.4]
  input  [31:0] io_b, // @[:@22977.4]
  input         io_flow, // @[:@22977.4]
  output [31:0] io_result // @[:@22977.4]
);
  wire  x395_mul_clock; // @[BigIPZynq.scala 63:21:@22992.4]
  wire  x395_mul_io_flow; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] x395_mul_io_a; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] x395_mul_io_b; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] x395_mul_io_out; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@23000.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@23000.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@22984.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@22986.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@22988.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@22990.4]
  Multiplier_9 x395_mul ( // @[BigIPZynq.scala 63:21:@22992.4]
    .clock(x395_mul_clock),
    .io_flow(x395_mul_io_flow),
    .io_a(x395_mul_io_a),
    .io_b(x395_mul_io_b),
    .io_out(x395_mul_io_out)
  );
  fix2fixBox_118 fix2fixBox ( // @[Math.scala 253:30:@23000.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@22984.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@22986.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@22988.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@22990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@23008.4]
  assign x395_mul_clock = clock; // @[:@22993.4]
  assign x395_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@22997.4]
  assign x395_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@22995.4]
  assign x395_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@22996.4]
  assign fix2fixBox_io_a = x395_mul_io_out; // @[Math.scala 254:23:@23003.4]
endmodule
module fix2fixBox_119( // @[:@23010.2]
  input  [31:0] io_a, // @[:@23013.4]
  output [31:0] io_b // @[:@23013.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@23025.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@23025.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@23028.4]
endmodule
module x396( // @[:@23030.2]
  input  [31:0] io_b, // @[:@23033.4]
  output [31:0] io_result // @[:@23033.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@23038.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@23038.4]
  fix2fixBox_119 fix2fixBox ( // @[BigIPZynq.scala 219:30:@23038.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@23046.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@23041.4]
endmodule
module RetimeWrapper_253( // @[:@23060.2]
  input         clock, // @[:@23061.4]
  input         reset, // @[:@23062.4]
  input         io_flow, // @[:@23063.4]
  input  [31:0] io_in, // @[:@23063.4]
  output [31:0] io_out // @[:@23063.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23065.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23065.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23065.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23065.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23065.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23065.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@23065.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23078.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23077.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@23076.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23075.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23074.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23072.4]
endmodule
module x397_sub( // @[:@23211.2]
  input         clock, // @[:@23212.4]
  input         reset, // @[:@23213.4]
  input  [31:0] io_a, // @[:@23214.4]
  input  [31:0] io_b, // @[:@23214.4]
  input         io_flow, // @[:@23214.4]
  output [31:0] io_result // @[:@23214.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@23222.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@23222.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@23229.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@23229.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@23240.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@23240.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@23240.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@23240.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@23240.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@23227.4 Math.scala 724:14:@23228.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@23234.4 Math.scala 724:14:@23235.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@23236.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@23237.4]
  __56 _ ( // @[Math.scala 720:24:@23222.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __56 __1 ( // @[Math.scala 720:24:@23229.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@23240.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@23227.4 Math.scala 724:14:@23228.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@23234.4 Math.scala 724:14:@23235.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@23236.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@23237.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@23248.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@23225.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@23232.4]
  assign fix2fixBox_clock = clock; // @[:@23241.4]
  assign fix2fixBox_reset = reset; // @[:@23242.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@23243.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@23246.4]
endmodule
module RetimeWrapper_259( // @[:@23684.2]
  input         clock, // @[:@23685.4]
  input         reset, // @[:@23686.4]
  input         io_flow, // @[:@23687.4]
  input  [31:0] io_in, // @[:@23687.4]
  output [31:0] io_out // @[:@23687.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23689.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23689.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23689.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23689.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23689.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23689.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@23689.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23702.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23701.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@23700.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23699.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23698.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23696.4]
endmodule
module RetimeWrapper_278( // @[:@26916.2]
  input         clock, // @[:@26917.4]
  input         reset, // @[:@26918.4]
  input         io_flow, // @[:@26919.4]
  input  [63:0] io_in, // @[:@26919.4]
  output [63:0] io_out // @[:@26919.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26921.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26921.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26921.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26921.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26921.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26921.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26921.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26934.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26933.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@26932.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26931.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26930.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26928.4]
endmodule
module x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@27032.2]
  input          clock, // @[:@27033.4]
  input          reset, // @[:@27034.4]
  output         io_in_x241_TREADY, // @[:@27035.4]
  input  [255:0] io_in_x241_TDATA, // @[:@27035.4]
  input  [7:0]   io_in_x241_TID, // @[:@27035.4]
  input  [7:0]   io_in_x241_TDEST, // @[:@27035.4]
  output         io_in_x242_TVALID, // @[:@27035.4]
  input          io_in_x242_TREADY, // @[:@27035.4]
  output [255:0] io_in_x242_TDATA, // @[:@27035.4]
  input          io_sigsIn_backpressure, // @[:@27035.4]
  input          io_sigsIn_datapathEn, // @[:@27035.4]
  input          io_sigsIn_break, // @[:@27035.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@27035.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@27035.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@27035.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@27035.4]
  input          io_rr // @[:@27035.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@27049.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@27049.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@27061.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@27061.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@27084.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@27084.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@27084.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@27084.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@27084.4]
  wire  x278_lb_0_clock; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_reset; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_11_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_11_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_11_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_11_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_11_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_11_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_10_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_10_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_10_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_10_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_10_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_10_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_9_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_9_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_9_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_9_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_9_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_9_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_8_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_8_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_8_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_8_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_8_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_8_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_7_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_7_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_7_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_7_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_7_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_7_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_6_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_6_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_6_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_6_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_6_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_6_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_5_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_5_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_5_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_5_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_5_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_5_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_4_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_4_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_4_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_4_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_4_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_4_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_3_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_3_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_3_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_3_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_3_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_3_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_2_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_2_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_2_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_2_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_2_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_2_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_1_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_1_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_1_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_1_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_1_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_1_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_0_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_rPort_0_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_rPort_0_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_0_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_rPort_0_backpressure; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_rPort_0_output_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_wPort_1_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_wPort_1_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_wPort_1_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_wPort_1_data_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_wPort_1_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_wPort_0_banks_1; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [2:0] x278_lb_0_io_wPort_0_banks_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [8:0] x278_lb_0_io_wPort_0_ofs_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire [31:0] x278_lb_0_io_wPort_0_data_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x278_lb_0_io_wPort_0_en_0; // @[m_x278_lb_0.scala 39:17:@27094.4]
  wire  x504_sub_1_clock; // @[Math.scala 191:24:@27257.4]
  wire  x504_sub_1_reset; // @[Math.scala 191:24:@27257.4]
  wire [31:0] x504_sub_1_io_a; // @[Math.scala 191:24:@27257.4]
  wire [31:0] x504_sub_1_io_b; // @[Math.scala 191:24:@27257.4]
  wire  x504_sub_1_io_flow; // @[Math.scala 191:24:@27257.4]
  wire [31:0] x504_sub_1_io_result; // @[Math.scala 191:24:@27257.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27284.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27284.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27284.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@27284.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@27284.4]
  wire  x287_sum_1_clock; // @[Math.scala 150:24:@27293.4]
  wire  x287_sum_1_reset; // @[Math.scala 150:24:@27293.4]
  wire [31:0] x287_sum_1_io_a; // @[Math.scala 150:24:@27293.4]
  wire [31:0] x287_sum_1_io_b; // @[Math.scala 150:24:@27293.4]
  wire  x287_sum_1_io_flow; // @[Math.scala 150:24:@27293.4]
  wire [31:0] x287_sum_1_io_result; // @[Math.scala 150:24:@27293.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@27303.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@27303.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@27303.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@27303.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@27303.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@27312.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@27312.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@27312.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@27312.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@27312.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@27321.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@27321.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@27321.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@27321.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@27321.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@27330.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@27330.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@27330.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@27330.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@27330.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@27339.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@27339.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@27339.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@27339.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@27339.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@27348.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@27348.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@27348.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@27348.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@27348.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@27359.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@27359.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@27359.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@27359.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@27359.4]
  wire  x289_rdcol_1_clock; // @[Math.scala 150:24:@27382.4]
  wire  x289_rdcol_1_reset; // @[Math.scala 150:24:@27382.4]
  wire [31:0] x289_rdcol_1_io_a; // @[Math.scala 150:24:@27382.4]
  wire [31:0] x289_rdcol_1_io_b; // @[Math.scala 150:24:@27382.4]
  wire  x289_rdcol_1_io_flow; // @[Math.scala 150:24:@27382.4]
  wire [31:0] x289_rdcol_1_io_result; // @[Math.scala 150:24:@27382.4]
  wire  x293_sum_1_clock; // @[Math.scala 150:24:@27422.4]
  wire  x293_sum_1_reset; // @[Math.scala 150:24:@27422.4]
  wire [31:0] x293_sum_1_io_a; // @[Math.scala 150:24:@27422.4]
  wire [31:0] x293_sum_1_io_b; // @[Math.scala 150:24:@27422.4]
  wire  x293_sum_1_io_flow; // @[Math.scala 150:24:@27422.4]
  wire [31:0] x293_sum_1_io_result; // @[Math.scala 150:24:@27422.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@27432.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@27432.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@27432.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@27432.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@27432.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@27441.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@27441.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@27441.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@27441.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@27441.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@27450.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@27450.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@27450.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@27450.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@27450.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@27461.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@27461.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@27461.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@27461.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@27461.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@27482.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@27482.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@27482.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@27482.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@27482.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@27498.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@27498.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@27498.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@27498.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@27498.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@27529.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@27529.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@27529.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@27529.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@27529.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@27538.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@27538.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@27556.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@27556.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@27556.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@27556.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@27556.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@27574.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@27574.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@27574.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@27574.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@27574.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@27586.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@27586.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@27586.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@27586.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@27586.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@27607.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@27607.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@27607.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@27607.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@27607.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@27631.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@27631.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@27631.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@27631.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@27631.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@27640.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@27640.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@27640.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@27640.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@27640.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@27649.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@27649.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@27649.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@27649.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@27649.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@27661.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@27661.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@27661.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@27661.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@27661.4]
  wire  x307_rdcol_1_clock; // @[Math.scala 150:24:@27684.4]
  wire  x307_rdcol_1_reset; // @[Math.scala 150:24:@27684.4]
  wire [31:0] x307_rdcol_1_io_a; // @[Math.scala 150:24:@27684.4]
  wire [31:0] x307_rdcol_1_io_b; // @[Math.scala 150:24:@27684.4]
  wire  x307_rdcol_1_io_flow; // @[Math.scala 150:24:@27684.4]
  wire [31:0] x307_rdcol_1_io_result; // @[Math.scala 150:24:@27684.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@27735.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@27735.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@27735.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@27735.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@27735.4]
  wire  x313_sum_1_clock; // @[Math.scala 150:24:@27744.4]
  wire  x313_sum_1_reset; // @[Math.scala 150:24:@27744.4]
  wire [31:0] x313_sum_1_io_a; // @[Math.scala 150:24:@27744.4]
  wire [31:0] x313_sum_1_io_b; // @[Math.scala 150:24:@27744.4]
  wire  x313_sum_1_io_flow; // @[Math.scala 150:24:@27744.4]
  wire [31:0] x313_sum_1_io_result; // @[Math.scala 150:24:@27744.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@27754.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@27754.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@27754.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@27754.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@27754.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@27763.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@27763.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@27763.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@27763.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@27763.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@27772.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@27772.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@27772.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@27772.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@27772.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@27784.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@27784.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@27784.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@27784.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@27784.4]
  wire  x316_rdcol_1_clock; // @[Math.scala 150:24:@27807.4]
  wire  x316_rdcol_1_reset; // @[Math.scala 150:24:@27807.4]
  wire [31:0] x316_rdcol_1_io_a; // @[Math.scala 150:24:@27807.4]
  wire [31:0] x316_rdcol_1_io_b; // @[Math.scala 150:24:@27807.4]
  wire  x316_rdcol_1_io_flow; // @[Math.scala 150:24:@27807.4]
  wire [31:0] x316_rdcol_1_io_result; // @[Math.scala 150:24:@27807.4]
  wire  x322_sum_1_clock; // @[Math.scala 150:24:@27858.4]
  wire  x322_sum_1_reset; // @[Math.scala 150:24:@27858.4]
  wire [31:0] x322_sum_1_io_a; // @[Math.scala 150:24:@27858.4]
  wire [31:0] x322_sum_1_io_b; // @[Math.scala 150:24:@27858.4]
  wire  x322_sum_1_io_flow; // @[Math.scala 150:24:@27858.4]
  wire [31:0] x322_sum_1_io_result; // @[Math.scala 150:24:@27858.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@27868.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@27868.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@27868.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@27868.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@27868.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@27877.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@27877.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@27877.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@27877.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@27877.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@27886.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@27886.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@27886.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@27886.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@27886.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@27898.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@27898.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@27898.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@27898.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@27898.4]
  wire  x325_rdrow_1_clock; // @[Math.scala 191:24:@27921.4]
  wire  x325_rdrow_1_reset; // @[Math.scala 191:24:@27921.4]
  wire [31:0] x325_rdrow_1_io_a; // @[Math.scala 191:24:@27921.4]
  wire [31:0] x325_rdrow_1_io_b; // @[Math.scala 191:24:@27921.4]
  wire  x325_rdrow_1_io_flow; // @[Math.scala 191:24:@27921.4]
  wire [31:0] x325_rdrow_1_io_result; // @[Math.scala 191:24:@27921.4]
  wire  x512_sub_1_clock; // @[Math.scala 191:24:@27993.4]
  wire  x512_sub_1_reset; // @[Math.scala 191:24:@27993.4]
  wire [31:0] x512_sub_1_io_a; // @[Math.scala 191:24:@27993.4]
  wire [31:0] x512_sub_1_io_b; // @[Math.scala 191:24:@27993.4]
  wire  x512_sub_1_io_flow; // @[Math.scala 191:24:@27993.4]
  wire [31:0] x512_sub_1_io_result; // @[Math.scala 191:24:@27993.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@28003.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@28003.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@28003.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@28003.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@28003.4]
  wire  x333_sum_1_clock; // @[Math.scala 150:24:@28012.4]
  wire  x333_sum_1_reset; // @[Math.scala 150:24:@28012.4]
  wire [31:0] x333_sum_1_io_a; // @[Math.scala 150:24:@28012.4]
  wire [31:0] x333_sum_1_io_b; // @[Math.scala 150:24:@28012.4]
  wire  x333_sum_1_io_flow; // @[Math.scala 150:24:@28012.4]
  wire [31:0] x333_sum_1_io_result; // @[Math.scala 150:24:@28012.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@28022.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@28022.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@28022.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@28022.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@28022.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@28031.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@28031.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@28031.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@28031.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@28031.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@28043.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@28043.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@28043.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@28043.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@28043.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@28064.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@28064.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@28064.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@28064.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@28064.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@28079.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@28079.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@28079.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@28079.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@28079.4]
  wire  x338_sum_1_clock; // @[Math.scala 150:24:@28090.4]
  wire  x338_sum_1_reset; // @[Math.scala 150:24:@28090.4]
  wire [31:0] x338_sum_1_io_a; // @[Math.scala 150:24:@28090.4]
  wire [31:0] x338_sum_1_io_b; // @[Math.scala 150:24:@28090.4]
  wire  x338_sum_1_io_flow; // @[Math.scala 150:24:@28090.4]
  wire [31:0] x338_sum_1_io_result; // @[Math.scala 150:24:@28090.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@28100.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@28100.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@28100.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@28100.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@28100.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@28112.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@28112.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@28112.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@28112.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@28112.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@28139.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@28139.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@28139.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@28139.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@28139.4]
  wire  x343_sum_1_clock; // @[Math.scala 150:24:@28148.4]
  wire  x343_sum_1_reset; // @[Math.scala 150:24:@28148.4]
  wire [31:0] x343_sum_1_io_a; // @[Math.scala 150:24:@28148.4]
  wire [31:0] x343_sum_1_io_b; // @[Math.scala 150:24:@28148.4]
  wire  x343_sum_1_io_flow; // @[Math.scala 150:24:@28148.4]
  wire [31:0] x343_sum_1_io_result; // @[Math.scala 150:24:@28148.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@28158.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@28158.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@28158.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@28158.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@28158.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@28170.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@28170.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@28170.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@28170.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@28170.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@28197.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@28197.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@28197.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@28197.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@28197.4]
  wire  x348_sum_1_clock; // @[Math.scala 150:24:@28206.4]
  wire  x348_sum_1_reset; // @[Math.scala 150:24:@28206.4]
  wire [31:0] x348_sum_1_io_a; // @[Math.scala 150:24:@28206.4]
  wire [31:0] x348_sum_1_io_b; // @[Math.scala 150:24:@28206.4]
  wire  x348_sum_1_io_flow; // @[Math.scala 150:24:@28206.4]
  wire [31:0] x348_sum_1_io_result; // @[Math.scala 150:24:@28206.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@28228.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@28228.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@28228.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@28228.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@28228.4]
  wire  x351_rdrow_1_clock; // @[Math.scala 191:24:@28251.4]
  wire  x351_rdrow_1_reset; // @[Math.scala 191:24:@28251.4]
  wire [31:0] x351_rdrow_1_io_a; // @[Math.scala 191:24:@28251.4]
  wire [31:0] x351_rdrow_1_io_b; // @[Math.scala 191:24:@28251.4]
  wire  x351_rdrow_1_io_flow; // @[Math.scala 191:24:@28251.4]
  wire [31:0] x351_rdrow_1_io_result; // @[Math.scala 191:24:@28251.4]
  wire  x517_sub_1_clock; // @[Math.scala 191:24:@28323.4]
  wire  x517_sub_1_reset; // @[Math.scala 191:24:@28323.4]
  wire [31:0] x517_sub_1_io_a; // @[Math.scala 191:24:@28323.4]
  wire [31:0] x517_sub_1_io_b; // @[Math.scala 191:24:@28323.4]
  wire  x517_sub_1_io_flow; // @[Math.scala 191:24:@28323.4]
  wire [31:0] x517_sub_1_io_result; // @[Math.scala 191:24:@28323.4]
  wire  x359_sum_1_clock; // @[Math.scala 150:24:@28333.4]
  wire  x359_sum_1_reset; // @[Math.scala 150:24:@28333.4]
  wire [31:0] x359_sum_1_io_a; // @[Math.scala 150:24:@28333.4]
  wire [31:0] x359_sum_1_io_b; // @[Math.scala 150:24:@28333.4]
  wire  x359_sum_1_io_flow; // @[Math.scala 150:24:@28333.4]
  wire [31:0] x359_sum_1_io_result; // @[Math.scala 150:24:@28333.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@28343.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@28343.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@28343.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@28343.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@28343.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@28352.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@28352.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@28352.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@28352.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@28352.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@28364.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@28364.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@28364.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@28364.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@28364.4]
  wire  x364_sum_1_clock; // @[Math.scala 150:24:@28391.4]
  wire  x364_sum_1_reset; // @[Math.scala 150:24:@28391.4]
  wire [31:0] x364_sum_1_io_a; // @[Math.scala 150:24:@28391.4]
  wire [31:0] x364_sum_1_io_b; // @[Math.scala 150:24:@28391.4]
  wire  x364_sum_1_io_flow; // @[Math.scala 150:24:@28391.4]
  wire [31:0] x364_sum_1_io_result; // @[Math.scala 150:24:@28391.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@28401.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@28401.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@28401.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@28401.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@28401.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@28413.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@28413.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@28413.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@28413.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@28413.4]
  wire  x369_sum_1_clock; // @[Math.scala 150:24:@28440.4]
  wire  x369_sum_1_reset; // @[Math.scala 150:24:@28440.4]
  wire [31:0] x369_sum_1_io_a; // @[Math.scala 150:24:@28440.4]
  wire [31:0] x369_sum_1_io_b; // @[Math.scala 150:24:@28440.4]
  wire  x369_sum_1_io_flow; // @[Math.scala 150:24:@28440.4]
  wire [31:0] x369_sum_1_io_result; // @[Math.scala 150:24:@28440.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@28450.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@28450.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@28450.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@28450.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@28450.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@28462.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@28462.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@28462.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@28462.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@28462.4]
  wire  x374_sum_1_clock; // @[Math.scala 150:24:@28491.4]
  wire  x374_sum_1_reset; // @[Math.scala 150:24:@28491.4]
  wire [31:0] x374_sum_1_io_a; // @[Math.scala 150:24:@28491.4]
  wire [31:0] x374_sum_1_io_b; // @[Math.scala 150:24:@28491.4]
  wire  x374_sum_1_io_flow; // @[Math.scala 150:24:@28491.4]
  wire [31:0] x374_sum_1_io_result; // @[Math.scala 150:24:@28491.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@28501.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@28501.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@28501.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@28501.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@28501.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@28513.4]
  wire  x377_1_clock; // @[Math.scala 262:24:@28536.4]
  wire [31:0] x377_1_io_a; // @[Math.scala 262:24:@28536.4]
  wire [31:0] x377_1_io_b; // @[Math.scala 262:24:@28536.4]
  wire  x377_1_io_flow; // @[Math.scala 262:24:@28536.4]
  wire [31:0] x377_1_io_result; // @[Math.scala 262:24:@28536.4]
  wire  x378_1_clock; // @[Math.scala 262:24:@28548.4]
  wire [31:0] x378_1_io_a; // @[Math.scala 262:24:@28548.4]
  wire [31:0] x378_1_io_b; // @[Math.scala 262:24:@28548.4]
  wire  x378_1_io_flow; // @[Math.scala 262:24:@28548.4]
  wire [31:0] x378_1_io_result; // @[Math.scala 262:24:@28548.4]
  wire  x379_1_clock; // @[Math.scala 262:24:@28560.4]
  wire [31:0] x379_1_io_a; // @[Math.scala 262:24:@28560.4]
  wire [31:0] x379_1_io_b; // @[Math.scala 262:24:@28560.4]
  wire  x379_1_io_flow; // @[Math.scala 262:24:@28560.4]
  wire [31:0] x379_1_io_result; // @[Math.scala 262:24:@28560.4]
  wire  x380_1_clock; // @[Math.scala 262:24:@28572.4]
  wire [31:0] x380_1_io_a; // @[Math.scala 262:24:@28572.4]
  wire [31:0] x380_1_io_b; // @[Math.scala 262:24:@28572.4]
  wire  x380_1_io_flow; // @[Math.scala 262:24:@28572.4]
  wire [31:0] x380_1_io_result; // @[Math.scala 262:24:@28572.4]
  wire  x381_1_clock; // @[Math.scala 262:24:@28584.4]
  wire [31:0] x381_1_io_a; // @[Math.scala 262:24:@28584.4]
  wire [31:0] x381_1_io_b; // @[Math.scala 262:24:@28584.4]
  wire  x381_1_io_flow; // @[Math.scala 262:24:@28584.4]
  wire [31:0] x381_1_io_result; // @[Math.scala 262:24:@28584.4]
  wire  x382_1_clock; // @[Math.scala 262:24:@28596.4]
  wire [31:0] x382_1_io_a; // @[Math.scala 262:24:@28596.4]
  wire [31:0] x382_1_io_b; // @[Math.scala 262:24:@28596.4]
  wire  x382_1_io_flow; // @[Math.scala 262:24:@28596.4]
  wire [31:0] x382_1_io_result; // @[Math.scala 262:24:@28596.4]
  wire  x383_1_clock; // @[Math.scala 262:24:@28608.4]
  wire [31:0] x383_1_io_a; // @[Math.scala 262:24:@28608.4]
  wire [31:0] x383_1_io_b; // @[Math.scala 262:24:@28608.4]
  wire  x383_1_io_flow; // @[Math.scala 262:24:@28608.4]
  wire [31:0] x383_1_io_result; // @[Math.scala 262:24:@28608.4]
  wire  x384_1_clock; // @[Math.scala 262:24:@28620.4]
  wire [31:0] x384_1_io_a; // @[Math.scala 262:24:@28620.4]
  wire [31:0] x384_1_io_b; // @[Math.scala 262:24:@28620.4]
  wire  x384_1_io_flow; // @[Math.scala 262:24:@28620.4]
  wire [31:0] x384_1_io_result; // @[Math.scala 262:24:@28620.4]
  wire  x385_1_clock; // @[Math.scala 262:24:@28632.4]
  wire [31:0] x385_1_io_a; // @[Math.scala 262:24:@28632.4]
  wire [31:0] x385_1_io_b; // @[Math.scala 262:24:@28632.4]
  wire  x385_1_io_flow; // @[Math.scala 262:24:@28632.4]
  wire [31:0] x385_1_io_result; // @[Math.scala 262:24:@28632.4]
  wire  x386_x13_1_clock; // @[Math.scala 150:24:@28642.4]
  wire  x386_x13_1_reset; // @[Math.scala 150:24:@28642.4]
  wire [31:0] x386_x13_1_io_a; // @[Math.scala 150:24:@28642.4]
  wire [31:0] x386_x13_1_io_b; // @[Math.scala 150:24:@28642.4]
  wire  x386_x13_1_io_flow; // @[Math.scala 150:24:@28642.4]
  wire [31:0] x386_x13_1_io_result; // @[Math.scala 150:24:@28642.4]
  wire  x387_x14_1_clock; // @[Math.scala 150:24:@28652.4]
  wire  x387_x14_1_reset; // @[Math.scala 150:24:@28652.4]
  wire [31:0] x387_x14_1_io_a; // @[Math.scala 150:24:@28652.4]
  wire [31:0] x387_x14_1_io_b; // @[Math.scala 150:24:@28652.4]
  wire  x387_x14_1_io_flow; // @[Math.scala 150:24:@28652.4]
  wire [31:0] x387_x14_1_io_result; // @[Math.scala 150:24:@28652.4]
  wire  x388_x13_1_clock; // @[Math.scala 150:24:@28662.4]
  wire  x388_x13_1_reset; // @[Math.scala 150:24:@28662.4]
  wire [31:0] x388_x13_1_io_a; // @[Math.scala 150:24:@28662.4]
  wire [31:0] x388_x13_1_io_b; // @[Math.scala 150:24:@28662.4]
  wire  x388_x13_1_io_flow; // @[Math.scala 150:24:@28662.4]
  wire [31:0] x388_x13_1_io_result; // @[Math.scala 150:24:@28662.4]
  wire  x389_x14_1_clock; // @[Math.scala 150:24:@28672.4]
  wire  x389_x14_1_reset; // @[Math.scala 150:24:@28672.4]
  wire [31:0] x389_x14_1_io_a; // @[Math.scala 150:24:@28672.4]
  wire [31:0] x389_x14_1_io_b; // @[Math.scala 150:24:@28672.4]
  wire  x389_x14_1_io_flow; // @[Math.scala 150:24:@28672.4]
  wire [31:0] x389_x14_1_io_result; // @[Math.scala 150:24:@28672.4]
  wire  x390_x13_1_clock; // @[Math.scala 150:24:@28682.4]
  wire  x390_x13_1_reset; // @[Math.scala 150:24:@28682.4]
  wire [31:0] x390_x13_1_io_a; // @[Math.scala 150:24:@28682.4]
  wire [31:0] x390_x13_1_io_b; // @[Math.scala 150:24:@28682.4]
  wire  x390_x13_1_io_flow; // @[Math.scala 150:24:@28682.4]
  wire [31:0] x390_x13_1_io_result; // @[Math.scala 150:24:@28682.4]
  wire  x391_x14_1_clock; // @[Math.scala 150:24:@28692.4]
  wire  x391_x14_1_reset; // @[Math.scala 150:24:@28692.4]
  wire [31:0] x391_x14_1_io_a; // @[Math.scala 150:24:@28692.4]
  wire [31:0] x391_x14_1_io_b; // @[Math.scala 150:24:@28692.4]
  wire  x391_x14_1_io_flow; // @[Math.scala 150:24:@28692.4]
  wire [31:0] x391_x14_1_io_result; // @[Math.scala 150:24:@28692.4]
  wire  x392_x13_1_clock; // @[Math.scala 150:24:@28702.4]
  wire  x392_x13_1_reset; // @[Math.scala 150:24:@28702.4]
  wire [31:0] x392_x13_1_io_a; // @[Math.scala 150:24:@28702.4]
  wire [31:0] x392_x13_1_io_b; // @[Math.scala 150:24:@28702.4]
  wire  x392_x13_1_io_flow; // @[Math.scala 150:24:@28702.4]
  wire [31:0] x392_x13_1_io_result; // @[Math.scala 150:24:@28702.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@28712.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@28712.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@28712.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@28712.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@28712.4]
  wire  x393_sum_1_clock; // @[Math.scala 150:24:@28721.4]
  wire  x393_sum_1_reset; // @[Math.scala 150:24:@28721.4]
  wire [31:0] x393_sum_1_io_a; // @[Math.scala 150:24:@28721.4]
  wire [31:0] x393_sum_1_io_b; // @[Math.scala 150:24:@28721.4]
  wire  x393_sum_1_io_flow; // @[Math.scala 150:24:@28721.4]
  wire [31:0] x393_sum_1_io_result; // @[Math.scala 150:24:@28721.4]
  wire [31:0] x394_1_io_b; // @[Math.scala 720:24:@28731.4]
  wire [31:0] x394_1_io_result; // @[Math.scala 720:24:@28731.4]
  wire  x395_mul_1_clock; // @[Math.scala 262:24:@28742.4]
  wire [31:0] x395_mul_1_io_a; // @[Math.scala 262:24:@28742.4]
  wire [31:0] x395_mul_1_io_b; // @[Math.scala 262:24:@28742.4]
  wire  x395_mul_1_io_flow; // @[Math.scala 262:24:@28742.4]
  wire [31:0] x395_mul_1_io_result; // @[Math.scala 262:24:@28742.4]
  wire [31:0] x396_1_io_b; // @[Math.scala 720:24:@28752.4]
  wire [31:0] x396_1_io_result; // @[Math.scala 720:24:@28752.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@28761.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@28761.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@28761.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@28761.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@28761.4]
  wire  x397_sub_1_clock; // @[Math.scala 191:24:@28770.4]
  wire  x397_sub_1_reset; // @[Math.scala 191:24:@28770.4]
  wire [31:0] x397_sub_1_io_a; // @[Math.scala 191:24:@28770.4]
  wire [31:0] x397_sub_1_io_b; // @[Math.scala 191:24:@28770.4]
  wire  x397_sub_1_io_flow; // @[Math.scala 191:24:@28770.4]
  wire [31:0] x397_sub_1_io_result; // @[Math.scala 191:24:@28770.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@28783.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@28783.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@28783.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@28783.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@28783.4]
  wire  x399_sub_1_clock; // @[Math.scala 191:24:@28792.4]
  wire  x399_sub_1_reset; // @[Math.scala 191:24:@28792.4]
  wire [31:0] x399_sub_1_io_a; // @[Math.scala 191:24:@28792.4]
  wire [31:0] x399_sub_1_io_b; // @[Math.scala 191:24:@28792.4]
  wire  x399_sub_1_io_flow; // @[Math.scala 191:24:@28792.4]
  wire [31:0] x399_sub_1_io_result; // @[Math.scala 191:24:@28792.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@28817.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@28817.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@28817.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@28817.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@28817.4]
  wire [31:0] x403_1_io_b; // @[Math.scala 720:24:@28831.4]
  wire [31:0] x403_1_io_result; // @[Math.scala 720:24:@28831.4]
  wire  x404_mul_1_clock; // @[Math.scala 262:24:@28842.4]
  wire [31:0] x404_mul_1_io_a; // @[Math.scala 262:24:@28842.4]
  wire [31:0] x404_mul_1_io_b; // @[Math.scala 262:24:@28842.4]
  wire  x404_mul_1_io_flow; // @[Math.scala 262:24:@28842.4]
  wire [31:0] x404_mul_1_io_result; // @[Math.scala 262:24:@28842.4]
  wire [31:0] x405_1_io_b; // @[Math.scala 720:24:@28852.4]
  wire [31:0] x405_1_io_result; // @[Math.scala 720:24:@28852.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@28861.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@28861.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@28861.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@28861.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@28861.4]
  wire  x406_sum_1_clock; // @[Math.scala 150:24:@28870.4]
  wire  x406_sum_1_reset; // @[Math.scala 150:24:@28870.4]
  wire [31:0] x406_sum_1_io_a; // @[Math.scala 150:24:@28870.4]
  wire [31:0] x406_sum_1_io_b; // @[Math.scala 150:24:@28870.4]
  wire  x406_sum_1_io_flow; // @[Math.scala 150:24:@28870.4]
  wire [31:0] x406_sum_1_io_result; // @[Math.scala 150:24:@28870.4]
  wire  x407_1_clock; // @[Math.scala 262:24:@28882.4]
  wire [31:0] x407_1_io_a; // @[Math.scala 262:24:@28882.4]
  wire [31:0] x407_1_io_b; // @[Math.scala 262:24:@28882.4]
  wire  x407_1_io_flow; // @[Math.scala 262:24:@28882.4]
  wire [31:0] x407_1_io_result; // @[Math.scala 262:24:@28882.4]
  wire  x408_1_clock; // @[Math.scala 262:24:@28894.4]
  wire [31:0] x408_1_io_a; // @[Math.scala 262:24:@28894.4]
  wire [31:0] x408_1_io_b; // @[Math.scala 262:24:@28894.4]
  wire  x408_1_io_flow; // @[Math.scala 262:24:@28894.4]
  wire [31:0] x408_1_io_result; // @[Math.scala 262:24:@28894.4]
  wire  x409_1_clock; // @[Math.scala 262:24:@28906.4]
  wire [31:0] x409_1_io_a; // @[Math.scala 262:24:@28906.4]
  wire [31:0] x409_1_io_b; // @[Math.scala 262:24:@28906.4]
  wire  x409_1_io_flow; // @[Math.scala 262:24:@28906.4]
  wire [31:0] x409_1_io_result; // @[Math.scala 262:24:@28906.4]
  wire  x410_1_clock; // @[Math.scala 262:24:@28918.4]
  wire [31:0] x410_1_io_a; // @[Math.scala 262:24:@28918.4]
  wire [31:0] x410_1_io_b; // @[Math.scala 262:24:@28918.4]
  wire  x410_1_io_flow; // @[Math.scala 262:24:@28918.4]
  wire [31:0] x410_1_io_result; // @[Math.scala 262:24:@28918.4]
  wire  x411_1_clock; // @[Math.scala 262:24:@28930.4]
  wire [31:0] x411_1_io_a; // @[Math.scala 262:24:@28930.4]
  wire [31:0] x411_1_io_b; // @[Math.scala 262:24:@28930.4]
  wire  x411_1_io_flow; // @[Math.scala 262:24:@28930.4]
  wire [31:0] x411_1_io_result; // @[Math.scala 262:24:@28930.4]
  wire  x412_1_clock; // @[Math.scala 262:24:@28942.4]
  wire [31:0] x412_1_io_a; // @[Math.scala 262:24:@28942.4]
  wire [31:0] x412_1_io_b; // @[Math.scala 262:24:@28942.4]
  wire  x412_1_io_flow; // @[Math.scala 262:24:@28942.4]
  wire [31:0] x412_1_io_result; // @[Math.scala 262:24:@28942.4]
  wire  x413_1_clock; // @[Math.scala 262:24:@28954.4]
  wire [31:0] x413_1_io_a; // @[Math.scala 262:24:@28954.4]
  wire [31:0] x413_1_io_b; // @[Math.scala 262:24:@28954.4]
  wire  x413_1_io_flow; // @[Math.scala 262:24:@28954.4]
  wire [31:0] x413_1_io_result; // @[Math.scala 262:24:@28954.4]
  wire  x414_1_clock; // @[Math.scala 262:24:@28966.4]
  wire [31:0] x414_1_io_a; // @[Math.scala 262:24:@28966.4]
  wire [31:0] x414_1_io_b; // @[Math.scala 262:24:@28966.4]
  wire  x414_1_io_flow; // @[Math.scala 262:24:@28966.4]
  wire [31:0] x414_1_io_result; // @[Math.scala 262:24:@28966.4]
  wire  x415_1_clock; // @[Math.scala 262:24:@28978.4]
  wire [31:0] x415_1_io_a; // @[Math.scala 262:24:@28978.4]
  wire [31:0] x415_1_io_b; // @[Math.scala 262:24:@28978.4]
  wire  x415_1_io_flow; // @[Math.scala 262:24:@28978.4]
  wire [31:0] x415_1_io_result; // @[Math.scala 262:24:@28978.4]
  wire  x416_x13_1_clock; // @[Math.scala 150:24:@28990.4]
  wire  x416_x13_1_reset; // @[Math.scala 150:24:@28990.4]
  wire [31:0] x416_x13_1_io_a; // @[Math.scala 150:24:@28990.4]
  wire [31:0] x416_x13_1_io_b; // @[Math.scala 150:24:@28990.4]
  wire  x416_x13_1_io_flow; // @[Math.scala 150:24:@28990.4]
  wire [31:0] x416_x13_1_io_result; // @[Math.scala 150:24:@28990.4]
  wire  x417_x14_1_clock; // @[Math.scala 150:24:@29000.4]
  wire  x417_x14_1_reset; // @[Math.scala 150:24:@29000.4]
  wire [31:0] x417_x14_1_io_a; // @[Math.scala 150:24:@29000.4]
  wire [31:0] x417_x14_1_io_b; // @[Math.scala 150:24:@29000.4]
  wire  x417_x14_1_io_flow; // @[Math.scala 150:24:@29000.4]
  wire [31:0] x417_x14_1_io_result; // @[Math.scala 150:24:@29000.4]
  wire  x418_x13_1_clock; // @[Math.scala 150:24:@29010.4]
  wire  x418_x13_1_reset; // @[Math.scala 150:24:@29010.4]
  wire [31:0] x418_x13_1_io_a; // @[Math.scala 150:24:@29010.4]
  wire [31:0] x418_x13_1_io_b; // @[Math.scala 150:24:@29010.4]
  wire  x418_x13_1_io_flow; // @[Math.scala 150:24:@29010.4]
  wire [31:0] x418_x13_1_io_result; // @[Math.scala 150:24:@29010.4]
  wire  x419_x14_1_clock; // @[Math.scala 150:24:@29020.4]
  wire  x419_x14_1_reset; // @[Math.scala 150:24:@29020.4]
  wire [31:0] x419_x14_1_io_a; // @[Math.scala 150:24:@29020.4]
  wire [31:0] x419_x14_1_io_b; // @[Math.scala 150:24:@29020.4]
  wire  x419_x14_1_io_flow; // @[Math.scala 150:24:@29020.4]
  wire [31:0] x419_x14_1_io_result; // @[Math.scala 150:24:@29020.4]
  wire  x420_x13_1_clock; // @[Math.scala 150:24:@29030.4]
  wire  x420_x13_1_reset; // @[Math.scala 150:24:@29030.4]
  wire [31:0] x420_x13_1_io_a; // @[Math.scala 150:24:@29030.4]
  wire [31:0] x420_x13_1_io_b; // @[Math.scala 150:24:@29030.4]
  wire  x420_x13_1_io_flow; // @[Math.scala 150:24:@29030.4]
  wire [31:0] x420_x13_1_io_result; // @[Math.scala 150:24:@29030.4]
  wire  x421_x14_1_clock; // @[Math.scala 150:24:@29040.4]
  wire  x421_x14_1_reset; // @[Math.scala 150:24:@29040.4]
  wire [31:0] x421_x14_1_io_a; // @[Math.scala 150:24:@29040.4]
  wire [31:0] x421_x14_1_io_b; // @[Math.scala 150:24:@29040.4]
  wire  x421_x14_1_io_flow; // @[Math.scala 150:24:@29040.4]
  wire [31:0] x421_x14_1_io_result; // @[Math.scala 150:24:@29040.4]
  wire  x422_x13_1_clock; // @[Math.scala 150:24:@29050.4]
  wire  x422_x13_1_reset; // @[Math.scala 150:24:@29050.4]
  wire [31:0] x422_x13_1_io_a; // @[Math.scala 150:24:@29050.4]
  wire [31:0] x422_x13_1_io_b; // @[Math.scala 150:24:@29050.4]
  wire  x422_x13_1_io_flow; // @[Math.scala 150:24:@29050.4]
  wire [31:0] x422_x13_1_io_result; // @[Math.scala 150:24:@29050.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@29060.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@29060.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@29060.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@29060.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@29060.4]
  wire  x423_sum_1_clock; // @[Math.scala 150:24:@29069.4]
  wire  x423_sum_1_reset; // @[Math.scala 150:24:@29069.4]
  wire [31:0] x423_sum_1_io_a; // @[Math.scala 150:24:@29069.4]
  wire [31:0] x423_sum_1_io_b; // @[Math.scala 150:24:@29069.4]
  wire  x423_sum_1_io_flow; // @[Math.scala 150:24:@29069.4]
  wire [31:0] x423_sum_1_io_result; // @[Math.scala 150:24:@29069.4]
  wire [31:0] x424_1_io_b; // @[Math.scala 720:24:@29079.4]
  wire [31:0] x424_1_io_result; // @[Math.scala 720:24:@29079.4]
  wire  x425_mul_1_clock; // @[Math.scala 262:24:@29090.4]
  wire [31:0] x425_mul_1_io_a; // @[Math.scala 262:24:@29090.4]
  wire [31:0] x425_mul_1_io_b; // @[Math.scala 262:24:@29090.4]
  wire  x425_mul_1_io_flow; // @[Math.scala 262:24:@29090.4]
  wire [31:0] x425_mul_1_io_result; // @[Math.scala 262:24:@29090.4]
  wire [31:0] x426_1_io_b; // @[Math.scala 720:24:@29100.4]
  wire [31:0] x426_1_io_result; // @[Math.scala 720:24:@29100.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@29109.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@29109.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@29109.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@29109.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@29109.4]
  wire  x427_sub_1_clock; // @[Math.scala 191:24:@29118.4]
  wire  x427_sub_1_reset; // @[Math.scala 191:24:@29118.4]
  wire [31:0] x427_sub_1_io_a; // @[Math.scala 191:24:@29118.4]
  wire [31:0] x427_sub_1_io_b; // @[Math.scala 191:24:@29118.4]
  wire  x427_sub_1_io_flow; // @[Math.scala 191:24:@29118.4]
  wire [31:0] x427_sub_1_io_result; // @[Math.scala 191:24:@29118.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@29131.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@29131.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@29131.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@29131.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@29131.4]
  wire  x429_sub_1_clock; // @[Math.scala 191:24:@29140.4]
  wire  x429_sub_1_reset; // @[Math.scala 191:24:@29140.4]
  wire [31:0] x429_sub_1_io_a; // @[Math.scala 191:24:@29140.4]
  wire [31:0] x429_sub_1_io_b; // @[Math.scala 191:24:@29140.4]
  wire  x429_sub_1_io_flow; // @[Math.scala 191:24:@29140.4]
  wire [31:0] x429_sub_1_io_result; // @[Math.scala 191:24:@29140.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@29153.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@29153.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@29153.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@29153.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@29153.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@29165.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@29165.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@29165.4]
  wire [31:0] RetimeWrapper_70_io_in; // @[package.scala 93:22:@29165.4]
  wire [31:0] RetimeWrapper_70_io_out; // @[package.scala 93:22:@29165.4]
  wire [31:0] x433_1_io_b; // @[Math.scala 720:24:@29179.4]
  wire [31:0] x433_1_io_result; // @[Math.scala 720:24:@29179.4]
  wire  x434_mul_1_clock; // @[Math.scala 262:24:@29190.4]
  wire [31:0] x434_mul_1_io_a; // @[Math.scala 262:24:@29190.4]
  wire [31:0] x434_mul_1_io_b; // @[Math.scala 262:24:@29190.4]
  wire  x434_mul_1_io_flow; // @[Math.scala 262:24:@29190.4]
  wire [31:0] x434_mul_1_io_result; // @[Math.scala 262:24:@29190.4]
  wire [31:0] x435_1_io_b; // @[Math.scala 720:24:@29200.4]
  wire [31:0] x435_1_io_result; // @[Math.scala 720:24:@29200.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@29209.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@29209.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@29209.4]
  wire [31:0] RetimeWrapper_71_io_in; // @[package.scala 93:22:@29209.4]
  wire [31:0] RetimeWrapper_71_io_out; // @[package.scala 93:22:@29209.4]
  wire  x436_sum_1_clock; // @[Math.scala 150:24:@29218.4]
  wire  x436_sum_1_reset; // @[Math.scala 150:24:@29218.4]
  wire [31:0] x436_sum_1_io_a; // @[Math.scala 150:24:@29218.4]
  wire [31:0] x436_sum_1_io_b; // @[Math.scala 150:24:@29218.4]
  wire  x436_sum_1_io_flow; // @[Math.scala 150:24:@29218.4]
  wire [31:0] x436_sum_1_io_result; // @[Math.scala 150:24:@29218.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@29234.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@29234.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@29234.4]
  wire [63:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@29234.4]
  wire [63:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@29234.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@29261.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@29261.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@29261.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@29261.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@29261.4]
  wire  b274; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 62:18:@27069.4]
  wire  b275; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 63:18:@27070.4]
  wire  _T_205; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 67:30:@27072.4]
  wire  _T_206; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 67:37:@27073.4]
  wire  _T_210; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 69:76:@27078.4]
  wire  _T_211; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 69:62:@27079.4]
  wire  _T_213; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 69:101:@27080.4]
  wire [63:0] x523_x276_D1_0_number; // @[package.scala 96:25:@27089.4 package.scala 96:25:@27090.4]
  wire [31:0] b272_number; // @[Math.scala 723:22:@27054.4 Math.scala 724:14:@27055.4]
  wire [31:0] _T_243; // @[Math.scala 406:49:@27198.4]
  wire [31:0] _T_245; // @[Math.scala 406:56:@27200.4]
  wire [31:0] _T_246; // @[Math.scala 406:56:@27201.4]
  wire [31:0] x499_number; // @[implicits.scala 133:21:@27202.4]
  wire [31:0] _T_256; // @[Math.scala 406:49:@27211.4]
  wire [31:0] _T_258; // @[Math.scala 406:56:@27213.4]
  wire [31:0] _T_259; // @[Math.scala 406:56:@27214.4]
  wire [31:0] b273_number; // @[Math.scala 723:22:@27066.4 Math.scala 724:14:@27067.4]
  wire [31:0] _T_268; // @[Math.scala 406:49:@27222.4]
  wire [31:0] _T_270; // @[Math.scala 406:56:@27224.4]
  wire [31:0] _T_271; // @[Math.scala 406:56:@27225.4]
  wire  _T_275; // @[FixedPoint.scala 50:25:@27231.4]
  wire [1:0] _T_279; // @[Bitwise.scala 72:12:@27233.4]
  wire [29:0] _T_280; // @[FixedPoint.scala 18:52:@27234.4]
  wire  _T_286; // @[Math.scala 451:55:@27236.4]
  wire [1:0] _T_287; // @[FixedPoint.scala 18:52:@27237.4]
  wire  _T_293; // @[Math.scala 451:110:@27239.4]
  wire  _T_294; // @[Math.scala 451:94:@27240.4]
  wire [31:0] _T_296; // @[Cat.scala 30:58:@27242.4]
  wire [31:0] x284_1_number; // @[Math.scala 454:20:@27243.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@27248.4]
  wire [40:0] _T_301; // @[Math.scala 461:32:@27248.4]
  wire [36:0] _GEN_1; // @[Math.scala 461:32:@27253.4]
  wire [36:0] _T_304; // @[Math.scala 461:32:@27253.4]
  wire  _T_310; // @[FixedPoint.scala 50:25:@27268.4]
  wire [1:0] _T_314; // @[Bitwise.scala 72:12:@27270.4]
  wire [29:0] _T_315; // @[FixedPoint.scala 18:52:@27271.4]
  wire  _T_321; // @[Math.scala 451:55:@27273.4]
  wire [1:0] _T_322; // @[FixedPoint.scala 18:52:@27274.4]
  wire  _T_328; // @[Math.scala 451:110:@27276.4]
  wire  _T_329; // @[Math.scala 451:94:@27277.4]
  wire [31:0] _T_331; // @[Cat.scala 30:58:@27279.4]
  wire  _T_359; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:101:@27356.4]
  wire  _T_363; // @[package.scala 96:25:@27364.4 package.scala 96:25:@27365.4]
  wire  _T_365; // @[implicits.scala 55:10:@27366.4]
  wire  _T_366; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:118:@27367.4]
  wire  _T_368; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:206:@27369.4]
  wire  _T_369; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:225:@27370.4]
  wire  x528_b274_D3; // @[package.scala 96:25:@27335.4 package.scala 96:25:@27336.4]
  wire  _T_370; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:251:@27371.4]
  wire  x526_b275_D3; // @[package.scala 96:25:@27317.4 package.scala 96:25:@27318.4]
  wire [31:0] x289_rdcol_number; // @[Math.scala 154:22:@27388.4 Math.scala 155:14:@27389.4]
  wire [31:0] _T_387; // @[Math.scala 406:49:@27397.4]
  wire [31:0] _T_389; // @[Math.scala 406:56:@27399.4]
  wire [31:0] _T_390; // @[Math.scala 406:56:@27400.4]
  wire  _T_394; // @[FixedPoint.scala 50:25:@27406.4]
  wire [1:0] _T_398; // @[Bitwise.scala 72:12:@27408.4]
  wire [29:0] _T_399; // @[FixedPoint.scala 18:52:@27409.4]
  wire  _T_405; // @[Math.scala 451:55:@27411.4]
  wire [1:0] _T_406; // @[FixedPoint.scala 18:52:@27412.4]
  wire  _T_412; // @[Math.scala 451:110:@27414.4]
  wire  _T_413; // @[Math.scala 451:94:@27415.4]
  wire [31:0] _T_415; // @[Cat.scala 30:58:@27417.4]
  wire  _T_435; // @[package.scala 96:25:@27466.4 package.scala 96:25:@27467.4]
  wire  _T_437; // @[implicits.scala 55:10:@27468.4]
  wire  _T_438; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:118:@27469.4]
  wire  _T_440; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:206:@27471.4]
  wire  _T_441; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:225:@27472.4]
  wire  _T_442; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:251:@27473.4]
  wire [31:0] x534_b272_D6_number; // @[package.scala 96:25:@27487.4 package.scala 96:25:@27488.4]
  wire [31:0] _T_452; // @[Math.scala 476:37:@27493.4]
  wire  x296; // @[Math.scala 476:44:@27495.4]
  wire [31:0] x535_x289_rdcol_D6_number; // @[package.scala 96:25:@27503.4 package.scala 96:25:@27504.4]
  wire [31:0] _T_463; // @[Math.scala 476:37:@27509.4]
  wire  x297; // @[Math.scala 476:44:@27511.4]
  wire  x536_x296_D1; // @[package.scala 96:25:@27519.4 package.scala 96:25:@27520.4]
  wire  x298; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 151:24:@27523.4]
  wire  _T_502; // @[package.scala 96:25:@27591.4 package.scala 96:25:@27592.4]
  wire  _T_504; // @[implicits.scala 55:10:@27593.4]
  wire  _T_505; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 170:146:@27594.4]
  wire  x541_x299_D2; // @[package.scala 96:25:@27570.4 package.scala 96:25:@27571.4]
  wire  _T_506; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 170:234:@27595.4]
  wire  x540_b274_D9; // @[package.scala 96:25:@27561.4 package.scala 96:25:@27562.4]
  wire  _T_507; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 170:242:@27596.4]
  wire  x539_b275_D9; // @[package.scala 96:25:@27552.4 package.scala 96:25:@27553.4]
  wire [31:0] x543_b273_D6_number; // @[package.scala 96:25:@27612.4 package.scala 96:25:@27613.4]
  wire [31:0] _T_520; // @[Math.scala 476:37:@27620.4]
  wire  x302; // @[Math.scala 476:44:@27622.4]
  wire  x303; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 186:59:@27625.4]
  wire  _T_547; // @[package.scala 96:25:@27666.4 package.scala 96:25:@27667.4]
  wire  _T_549; // @[implicits.scala 55:10:@27668.4]
  wire  _T_550; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 199:194:@27669.4]
  wire  x544_x304_D3; // @[package.scala 96:25:@27636.4 package.scala 96:25:@27637.4]
  wire  _T_551; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 199:282:@27670.4]
  wire  _T_552; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 199:290:@27671.4]
  wire [31:0] x307_rdcol_number; // @[Math.scala 154:22:@27690.4 Math.scala 155:14:@27691.4]
  wire [31:0] _T_567; // @[Math.scala 476:37:@27696.4]
  wire  x308; // @[Math.scala 476:44:@27698.4]
  wire  x309; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 207:59:@27701.4]
  wire [31:0] _T_583; // @[Math.scala 406:56:@27712.4]
  wire [31:0] _T_584; // @[Math.scala 406:56:@27713.4]
  wire  _T_588; // @[FixedPoint.scala 50:25:@27719.4]
  wire [1:0] _T_592; // @[Bitwise.scala 72:12:@27721.4]
  wire [29:0] _T_593; // @[FixedPoint.scala 18:52:@27722.4]
  wire  _T_599; // @[Math.scala 451:55:@27724.4]
  wire [1:0] _T_600; // @[FixedPoint.scala 18:52:@27725.4]
  wire  _T_606; // @[Math.scala 451:110:@27727.4]
  wire  _T_607; // @[Math.scala 451:94:@27728.4]
  wire [31:0] _T_609; // @[Cat.scala 30:58:@27730.4]
  wire  _T_638; // @[package.scala 96:25:@27789.4 package.scala 96:25:@27790.4]
  wire  _T_640; // @[implicits.scala 55:10:@27791.4]
  wire  _T_641; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 228:194:@27792.4]
  wire  x549_x310_D2; // @[package.scala 96:25:@27768.4 package.scala 96:25:@27769.4]
  wire  _T_642; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 228:282:@27793.4]
  wire  _T_643; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 228:290:@27794.4]
  wire [31:0] x316_rdcol_number; // @[Math.scala 154:22:@27813.4 Math.scala 155:14:@27814.4]
  wire [31:0] _T_658; // @[Math.scala 476:37:@27819.4]
  wire  x317; // @[Math.scala 476:44:@27821.4]
  wire  x318; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 236:59:@27824.4]
  wire [31:0] _T_674; // @[Math.scala 406:56:@27835.4]
  wire [31:0] _T_675; // @[Math.scala 406:56:@27836.4]
  wire  _T_679; // @[FixedPoint.scala 50:25:@27842.4]
  wire [1:0] _T_683; // @[Bitwise.scala 72:12:@27844.4]
  wire [29:0] _T_684; // @[FixedPoint.scala 18:52:@27845.4]
  wire  _T_690; // @[Math.scala 451:55:@27847.4]
  wire [1:0] _T_691; // @[FixedPoint.scala 18:52:@27848.4]
  wire  _T_697; // @[Math.scala 451:110:@27850.4]
  wire  _T_698; // @[Math.scala 451:94:@27851.4]
  wire [31:0] _T_700; // @[Cat.scala 30:58:@27853.4]
  wire  _T_726; // @[package.scala 96:25:@27903.4 package.scala 96:25:@27904.4]
  wire  _T_728; // @[implicits.scala 55:10:@27905.4]
  wire  _T_729; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 255:194:@27906.4]
  wire  x552_x319_D2; // @[package.scala 96:25:@27882.4 package.scala 96:25:@27883.4]
  wire  _T_730; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 255:282:@27907.4]
  wire  _T_731; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 255:290:@27908.4]
  wire [31:0] x325_rdrow_number; // @[Math.scala 195:22:@27927.4 Math.scala 196:14:@27928.4]
  wire [31:0] _T_748; // @[Math.scala 406:49:@27934.4]
  wire [31:0] _T_750; // @[Math.scala 406:56:@27936.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@27937.4]
  wire [31:0] x508_number; // @[implicits.scala 133:21:@27938.4]
  wire  x327; // @[Math.scala 476:44:@27946.4]
  wire  x328; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 265:24:@27949.4]
  wire [31:0] _T_772; // @[Math.scala 406:49:@27958.4]
  wire [31:0] _T_774; // @[Math.scala 406:56:@27960.4]
  wire [31:0] _T_775; // @[Math.scala 406:56:@27961.4]
  wire  _T_779; // @[FixedPoint.scala 50:25:@27967.4]
  wire [1:0] _T_783; // @[Bitwise.scala 72:12:@27969.4]
  wire [29:0] _T_784; // @[FixedPoint.scala 18:52:@27970.4]
  wire  _T_790; // @[Math.scala 451:55:@27972.4]
  wire [1:0] _T_791; // @[FixedPoint.scala 18:52:@27973.4]
  wire  _T_797; // @[Math.scala 451:110:@27975.4]
  wire  _T_798; // @[Math.scala 451:94:@27976.4]
  wire [31:0] _T_800; // @[Cat.scala 30:58:@27978.4]
  wire [31:0] x331_1_number; // @[Math.scala 454:20:@27979.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@27984.4]
  wire [40:0] _T_805; // @[Math.scala 461:32:@27984.4]
  wire [36:0] _GEN_3; // @[Math.scala 461:32:@27989.4]
  wire [36:0] _T_808; // @[Math.scala 461:32:@27989.4]
  wire  _T_835; // @[package.scala 96:25:@28048.4 package.scala 96:25:@28049.4]
  wire  _T_837; // @[implicits.scala 55:10:@28050.4]
  wire  _T_838; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 290:194:@28051.4]
  wire  x555_x329_D2; // @[package.scala 96:25:@28027.4 package.scala 96:25:@28028.4]
  wire  _T_839; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 290:282:@28052.4]
  wire  _T_840; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 290:290:@28053.4]
  wire  x557_x302_D1; // @[package.scala 96:25:@28069.4 package.scala 96:25:@28070.4]
  wire  x336; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 302:59:@28073.4]
  wire  _T_872; // @[package.scala 96:25:@28117.4 package.scala 96:25:@28118.4]
  wire  _T_874; // @[implicits.scala 55:10:@28119.4]
  wire  _T_875; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 317:194:@28120.4]
  wire  x559_x337_D2; // @[package.scala 96:25:@28105.4 package.scala 96:25:@28106.4]
  wire  _T_876; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 317:282:@28121.4]
  wire  _T_877; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 317:290:@28122.4]
  wire  x341; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 321:59:@28133.4]
  wire  _T_904; // @[package.scala 96:25:@28175.4 package.scala 96:25:@28176.4]
  wire  _T_906; // @[implicits.scala 55:10:@28177.4]
  wire  _T_907; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 334:194:@28178.4]
  wire  x561_x342_D2; // @[package.scala 96:25:@28163.4 package.scala 96:25:@28164.4]
  wire  _T_908; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 334:282:@28179.4]
  wire  _T_909; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 334:290:@28180.4]
  wire  x346; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 338:59:@28191.4]
  wire  _T_936; // @[package.scala 96:25:@28233.4 package.scala 96:25:@28234.4]
  wire  _T_938; // @[implicits.scala 55:10:@28235.4]
  wire  _T_939; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 351:194:@28236.4]
  wire  x563_x347_D2; // @[package.scala 96:25:@28221.4 package.scala 96:25:@28222.4]
  wire  _T_940; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 351:282:@28237.4]
  wire  _T_941; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 351:290:@28238.4]
  wire [31:0] x351_rdrow_number; // @[Math.scala 195:22:@28257.4 Math.scala 196:14:@28258.4]
  wire [31:0] _T_958; // @[Math.scala 406:49:@28264.4]
  wire [31:0] _T_960; // @[Math.scala 406:56:@28266.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@28267.4]
  wire [31:0] x513_number; // @[implicits.scala 133:21:@28268.4]
  wire  x353; // @[Math.scala 476:44:@28276.4]
  wire  x354; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 361:24:@28279.4]
  wire [31:0] _T_982; // @[Math.scala 406:49:@28288.4]
  wire [31:0] _T_984; // @[Math.scala 406:56:@28290.4]
  wire [31:0] _T_985; // @[Math.scala 406:56:@28291.4]
  wire  _T_989; // @[FixedPoint.scala 50:25:@28297.4]
  wire [1:0] _T_993; // @[Bitwise.scala 72:12:@28299.4]
  wire [29:0] _T_994; // @[FixedPoint.scala 18:52:@28300.4]
  wire  _T_1000; // @[Math.scala 451:55:@28302.4]
  wire [1:0] _T_1001; // @[FixedPoint.scala 18:52:@28303.4]
  wire  _T_1007; // @[Math.scala 451:110:@28305.4]
  wire  _T_1008; // @[Math.scala 451:94:@28306.4]
  wire [31:0] _T_1010; // @[Cat.scala 30:58:@28308.4]
  wire [31:0] x357_1_number; // @[Math.scala 454:20:@28309.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@28314.4]
  wire [40:0] _T_1015; // @[Math.scala 461:32:@28314.4]
  wire [36:0] _GEN_5; // @[Math.scala 461:32:@28319.4]
  wire [36:0] _T_1018; // @[Math.scala 461:32:@28319.4]
  wire  _T_1042; // @[package.scala 96:25:@28369.4 package.scala 96:25:@28370.4]
  wire  _T_1044; // @[implicits.scala 55:10:@28371.4]
  wire  _T_1045; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 384:194:@28372.4]
  wire  x565_x355_D2; // @[package.scala 96:25:@28357.4 package.scala 96:25:@28358.4]
  wire  _T_1046; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 384:282:@28373.4]
  wire  _T_1047; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 384:290:@28374.4]
  wire  x362; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 388:24:@28385.4]
  wire  _T_1071; // @[package.scala 96:25:@28418.4 package.scala 96:25:@28419.4]
  wire  _T_1073; // @[implicits.scala 55:10:@28420.4]
  wire  _T_1074; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 399:194:@28421.4]
  wire  x566_x363_D2; // @[package.scala 96:25:@28406.4 package.scala 96:25:@28407.4]
  wire  _T_1075; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 399:282:@28422.4]
  wire  _T_1076; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 399:290:@28423.4]
  wire  x367; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 403:24:@28434.4]
  wire  _T_1100; // @[package.scala 96:25:@28467.4 package.scala 96:25:@28468.4]
  wire  _T_1102; // @[implicits.scala 55:10:@28469.4]
  wire  _T_1103; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 414:194:@28470.4]
  wire  x567_x368_D2; // @[package.scala 96:25:@28455.4 package.scala 96:25:@28456.4]
  wire  _T_1104; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 414:282:@28471.4]
  wire  _T_1105; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 414:290:@28472.4]
  wire  x372; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 424:59:@28483.4]
  wire  _T_1131; // @[package.scala 96:25:@28518.4 package.scala 96:25:@28519.4]
  wire  _T_1133; // @[implicits.scala 55:10:@28520.4]
  wire  _T_1134; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 437:194:@28521.4]
  wire  x568_x373_D2; // @[package.scala 96:25:@28506.4 package.scala 96:25:@28507.4]
  wire  _T_1135; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 437:282:@28522.4]
  wire  _T_1136; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 437:290:@28523.4]
  wire [31:0] x397_sub_number; // @[Math.scala 195:22:@28776.4 Math.scala 196:14:@28777.4]
  wire [31:0] x399_sub_number; // @[Math.scala 195:22:@28798.4 Math.scala 196:14:@28799.4]
  wire  x398; // @[package.scala 96:25:@28788.4 package.scala 96:25:@28789.4]
  wire  x400; // @[package.scala 96:25:@28810.4 package.scala 96:25:@28811.4]
  wire  x401; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 493:24:@28814.4]
  wire [31:0] x571_x397_sub_D1_number; // @[package.scala 96:25:@28822.4 package.scala 96:25:@28823.4]
  wire [31:0] x427_sub_number; // @[Math.scala 195:22:@29124.4 Math.scala 196:14:@29125.4]
  wire [31:0] x429_sub_number; // @[Math.scala 195:22:@29146.4 Math.scala 196:14:@29147.4]
  wire  x428; // @[package.scala 96:25:@29136.4 package.scala 96:25:@29137.4]
  wire  x430; // @[package.scala 96:25:@29158.4 package.scala 96:25:@29159.4]
  wire  x431; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 569:24:@29162.4]
  wire [31:0] x575_x427_sub_D1_number; // @[package.scala 96:25:@29170.4 package.scala 96:25:@29171.4]
  wire [31:0] x406_sum_number; // @[Math.scala 154:22:@28876.4 Math.scala 155:14:@28877.4]
  wire [31:0] x436_sum_number; // @[Math.scala 154:22:@29224.4 Math.scala 155:14:@29225.4]
  wire  _T_1478; // @[package.scala 96:25:@29266.4 package.scala 96:25:@29267.4]
  wire  _T_1480; // @[implicits.scala 55:10:@29268.4]
  wire  x577_b274_D39; // @[package.scala 96:25:@29248.4 package.scala 96:25:@29249.4]
  wire  _T_1481; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 593:117:@29269.4]
  wire  x578_b275_D39; // @[package.scala 96:25:@29257.4 package.scala 96:25:@29258.4]
  wire  _T_1482; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 593:123:@29270.4]
  wire [31:0] x525_x500_D3_number; // @[package.scala 96:25:@27308.4 package.scala 96:25:@27309.4]
  wire [31:0] x529_x287_sum_D1_number; // @[package.scala 96:25:@27344.4 package.scala 96:25:@27345.4]
  wire [31:0] x530_x501_D3_number; // @[package.scala 96:25:@27353.4 package.scala 96:25:@27354.4]
  wire [31:0] x531_x293_sum_D1_number; // @[package.scala 96:25:@27437.4 package.scala 96:25:@27438.4]
  wire [31:0] x532_x505_D2_number; // @[package.scala 96:25:@27446.4 package.scala 96:25:@27447.4]
  wire [31:0] x537_x500_D9_number; // @[package.scala 96:25:@27534.4 package.scala 96:25:@27535.4]
  wire [31:0] x538_x293_sum_D7_number; // @[package.scala 96:25:@27543.4 package.scala 96:25:@27544.4]
  wire [31:0] x542_x505_D8_number; // @[package.scala 96:25:@27579.4 package.scala 96:25:@27580.4]
  wire [31:0] x545_x287_sum_D7_number; // @[package.scala 96:25:@27645.4 package.scala 96:25:@27646.4]
  wire [31:0] x546_x501_D9_number; // @[package.scala 96:25:@27654.4 package.scala 96:25:@27655.4]
  wire [31:0] x548_x313_sum_D1_number; // @[package.scala 96:25:@27759.4 package.scala 96:25:@27760.4]
  wire [31:0] x550_x506_D2_number; // @[package.scala 96:25:@27777.4 package.scala 96:25:@27778.4]
  wire [31:0] x551_x507_D2_number; // @[package.scala 96:25:@27873.4 package.scala 96:25:@27874.4]
  wire [31:0] x553_x322_sum_D1_number; // @[package.scala 96:25:@27891.4 package.scala 96:25:@27892.4]
  wire [31:0] x333_sum_number; // @[Math.scala 154:22:@28018.4 Math.scala 155:14:@28019.4]
  wire [31:0] x556_x509_D2_number; // @[package.scala 96:25:@28036.4 package.scala 96:25:@28037.4]
  wire [31:0] x338_sum_number; // @[Math.scala 154:22:@28096.4 Math.scala 155:14:@28097.4]
  wire [31:0] x343_sum_number; // @[Math.scala 154:22:@28154.4 Math.scala 155:14:@28155.4]
  wire [31:0] x348_sum_number; // @[Math.scala 154:22:@28212.4 Math.scala 155:14:@28213.4]
  wire [31:0] x359_sum_number; // @[Math.scala 154:22:@28339.4 Math.scala 155:14:@28340.4]
  wire [31:0] x564_x514_D2_number; // @[package.scala 96:25:@28348.4 package.scala 96:25:@28349.4]
  wire [31:0] x364_sum_number; // @[Math.scala 154:22:@28397.4 Math.scala 155:14:@28398.4]
  wire [31:0] x369_sum_number; // @[Math.scala 154:22:@28446.4 Math.scala 155:14:@28447.4]
  wire [31:0] x374_sum_number; // @[Math.scala 154:22:@28497.4 Math.scala 155:14:@28498.4]
  _ _ ( // @[Math.scala 720:24:@27049.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@27061.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@27084.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x278_lb_0 x278_lb_0 ( // @[m_x278_lb_0.scala 39:17:@27094.4]
    .clock(x278_lb_0_clock),
    .reset(x278_lb_0_reset),
    .io_rPort_11_banks_1(x278_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x278_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x278_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x278_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x278_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x278_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x278_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x278_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x278_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x278_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x278_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x278_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x278_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x278_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x278_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x278_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x278_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x278_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x278_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x278_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x278_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x278_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x278_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x278_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x278_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x278_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x278_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x278_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x278_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x278_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x278_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x278_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x278_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x278_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x278_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x278_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x278_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x278_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x278_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x278_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x278_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x278_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x278_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x278_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x278_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x278_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x278_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x278_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x278_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x278_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x278_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x278_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x278_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x278_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x278_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x278_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x278_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x278_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x278_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x278_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x278_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x278_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x278_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x278_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x278_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x278_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x278_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x278_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x278_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x278_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x278_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x278_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x278_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x278_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x278_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x278_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x278_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x278_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x278_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x278_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x278_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x278_lb_0_io_wPort_0_en_0)
  );
  x492_sub x504_sub_1 ( // @[Math.scala 191:24:@27257.4]
    .clock(x504_sub_1_clock),
    .reset(x504_sub_1_reset),
    .io_a(x504_sub_1_io_a),
    .io_b(x504_sub_1_io_b),
    .io_flow(x504_sub_1_io_flow),
    .io_result(x504_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@27284.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x255_sum x287_sum_1 ( // @[Math.scala 150:24:@27293.4]
    .clock(x287_sum_1_clock),
    .reset(x287_sum_1_reset),
    .io_a(x287_sum_1_io_a),
    .io_b(x287_sum_1_io_b),
    .io_flow(x287_sum_1_io_flow),
    .io_result(x287_sum_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_2 ( // @[package.scala 93:22:@27303.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_3 ( // @[package.scala 93:22:@27312.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_4 ( // @[package.scala 93:22:@27321.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_5 ( // @[package.scala 93:22:@27330.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_6 ( // @[package.scala 93:22:@27339.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_168 RetimeWrapper_7 ( // @[package.scala 93:22:@27348.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_8 ( // @[package.scala 93:22:@27359.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x255_sum x289_rdcol_1 ( // @[Math.scala 150:24:@27382.4]
    .clock(x289_rdcol_1_clock),
    .reset(x289_rdcol_1_reset),
    .io_a(x289_rdcol_1_io_a),
    .io_b(x289_rdcol_1_io_b),
    .io_flow(x289_rdcol_1_io_flow),
    .io_result(x289_rdcol_1_io_result)
  );
  x255_sum x293_sum_1 ( // @[Math.scala 150:24:@27422.4]
    .clock(x293_sum_1_clock),
    .reset(x293_sum_1_reset),
    .io_a(x293_sum_1_io_a),
    .io_b(x293_sum_1_io_b),
    .io_flow(x293_sum_1_io_flow),
    .io_result(x293_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_9 ( // @[package.scala 93:22:@27432.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_10 ( // @[package.scala 93:22:@27441.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_11 ( // @[package.scala 93:22:@27450.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_12 ( // @[package.scala 93:22:@27461.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_13 ( // @[package.scala 93:22:@27482.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_14 ( // @[package.scala 93:22:@27498.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@27514.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_184 RetimeWrapper_16 ( // @[package.scala 93:22:@27529.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_185 RetimeWrapper_17 ( // @[package.scala 93:22:@27538.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_18 ( // @[package.scala 93:22:@27547.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_19 ( // @[package.scala 93:22:@27556.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@27565.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_21 ( // @[package.scala 93:22:@27574.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_22 ( // @[package.scala 93:22:@27586.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_23 ( // @[package.scala 93:22:@27607.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_24 ( // @[package.scala 93:22:@27631.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_185 RetimeWrapper_25 ( // @[package.scala 93:22:@27640.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_184 RetimeWrapper_26 ( // @[package.scala 93:22:@27649.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_27 ( // @[package.scala 93:22:@27661.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x255_sum x307_rdcol_1 ( // @[Math.scala 150:24:@27684.4]
    .clock(x307_rdcol_1_clock),
    .reset(x307_rdcol_1_reset),
    .io_a(x307_rdcol_1_io_a),
    .io_b(x307_rdcol_1_io_b),
    .io_flow(x307_rdcol_1_io_flow),
    .io_result(x307_rdcol_1_io_result)
  );
  RetimeWrapper_181 RetimeWrapper_28 ( // @[package.scala 93:22:@27735.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x255_sum x313_sum_1 ( // @[Math.scala 150:24:@27744.4]
    .clock(x313_sum_1_clock),
    .reset(x313_sum_1_reset),
    .io_a(x313_sum_1_io_a),
    .io_b(x313_sum_1_io_b),
    .io_flow(x313_sum_1_io_flow),
    .io_result(x313_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_29 ( // @[package.scala 93:22:@27754.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@27763.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_31 ( // @[package.scala 93:22:@27772.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_32 ( // @[package.scala 93:22:@27784.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x255_sum x316_rdcol_1 ( // @[Math.scala 150:24:@27807.4]
    .clock(x316_rdcol_1_clock),
    .reset(x316_rdcol_1_reset),
    .io_a(x316_rdcol_1_io_a),
    .io_b(x316_rdcol_1_io_b),
    .io_flow(x316_rdcol_1_io_flow),
    .io_result(x316_rdcol_1_io_result)
  );
  x255_sum x322_sum_1 ( // @[Math.scala 150:24:@27858.4]
    .clock(x322_sum_1_clock),
    .reset(x322_sum_1_reset),
    .io_a(x322_sum_1_io_a),
    .io_b(x322_sum_1_io_b),
    .io_flow(x322_sum_1_io_flow),
    .io_result(x322_sum_1_io_result)
  );
  RetimeWrapper_170 RetimeWrapper_33 ( // @[package.scala 93:22:@27868.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@27877.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_35 ( // @[package.scala 93:22:@27886.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_36 ( // @[package.scala 93:22:@27898.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x492_sub x325_rdrow_1 ( // @[Math.scala 191:24:@27921.4]
    .clock(x325_rdrow_1_clock),
    .reset(x325_rdrow_1_reset),
    .io_a(x325_rdrow_1_io_a),
    .io_b(x325_rdrow_1_io_b),
    .io_flow(x325_rdrow_1_io_flow),
    .io_result(x325_rdrow_1_io_result)
  );
  x492_sub x512_sub_1 ( // @[Math.scala 191:24:@27993.4]
    .clock(x512_sub_1_clock),
    .reset(x512_sub_1_reset),
    .io_a(x512_sub_1_io_a),
    .io_b(x512_sub_1_io_b),
    .io_flow(x512_sub_1_io_flow),
    .io_result(x512_sub_1_io_result)
  );
  RetimeWrapper_185 RetimeWrapper_37 ( // @[package.scala 93:22:@28003.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x255_sum x333_sum_1 ( // @[Math.scala 150:24:@28012.4]
    .clock(x333_sum_1_clock),
    .reset(x333_sum_1_reset),
    .io_a(x333_sum_1_io_a),
    .io_b(x333_sum_1_io_b),
    .io_flow(x333_sum_1_io_flow),
    .io_result(x333_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@28022.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_39 ( // @[package.scala 93:22:@28031.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_40 ( // @[package.scala 93:22:@28043.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@28064.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_42 ( // @[package.scala 93:22:@28079.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  x255_sum x338_sum_1 ( // @[Math.scala 150:24:@28090.4]
    .clock(x338_sum_1_clock),
    .reset(x338_sum_1_reset),
    .io_a(x338_sum_1_io_a),
    .io_b(x338_sum_1_io_b),
    .io_flow(x338_sum_1_io_flow),
    .io_result(x338_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@28100.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_44 ( // @[package.scala 93:22:@28112.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_45 ( // @[package.scala 93:22:@28139.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x255_sum x343_sum_1 ( // @[Math.scala 150:24:@28148.4]
    .clock(x343_sum_1_clock),
    .reset(x343_sum_1_reset),
    .io_a(x343_sum_1_io_a),
    .io_b(x343_sum_1_io_b),
    .io_flow(x343_sum_1_io_flow),
    .io_result(x343_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@28158.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_47 ( // @[package.scala 93:22:@28170.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_48 ( // @[package.scala 93:22:@28197.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x255_sum x348_sum_1 ( // @[Math.scala 150:24:@28206.4]
    .clock(x348_sum_1_clock),
    .reset(x348_sum_1_reset),
    .io_a(x348_sum_1_io_a),
    .io_b(x348_sum_1_io_b),
    .io_flow(x348_sum_1_io_flow),
    .io_result(x348_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@28216.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_50 ( // @[package.scala 93:22:@28228.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x492_sub x351_rdrow_1 ( // @[Math.scala 191:24:@28251.4]
    .clock(x351_rdrow_1_clock),
    .reset(x351_rdrow_1_reset),
    .io_a(x351_rdrow_1_io_a),
    .io_b(x351_rdrow_1_io_b),
    .io_flow(x351_rdrow_1_io_flow),
    .io_result(x351_rdrow_1_io_result)
  );
  x492_sub x517_sub_1 ( // @[Math.scala 191:24:@28323.4]
    .clock(x517_sub_1_clock),
    .reset(x517_sub_1_reset),
    .io_a(x517_sub_1_io_a),
    .io_b(x517_sub_1_io_b),
    .io_flow(x517_sub_1_io_flow),
    .io_result(x517_sub_1_io_result)
  );
  x255_sum x359_sum_1 ( // @[Math.scala 150:24:@28333.4]
    .clock(x359_sum_1_clock),
    .reset(x359_sum_1_reset),
    .io_a(x359_sum_1_io_a),
    .io_b(x359_sum_1_io_b),
    .io_flow(x359_sum_1_io_flow),
    .io_result(x359_sum_1_io_result)
  );
  RetimeWrapper_170 RetimeWrapper_51 ( // @[package.scala 93:22:@28343.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@28352.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_53 ( // @[package.scala 93:22:@28364.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x255_sum x364_sum_1 ( // @[Math.scala 150:24:@28391.4]
    .clock(x364_sum_1_clock),
    .reset(x364_sum_1_reset),
    .io_a(x364_sum_1_io_a),
    .io_b(x364_sum_1_io_b),
    .io_flow(x364_sum_1_io_flow),
    .io_result(x364_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@28401.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_55 ( // @[package.scala 93:22:@28413.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x255_sum x369_sum_1 ( // @[Math.scala 150:24:@28440.4]
    .clock(x369_sum_1_clock),
    .reset(x369_sum_1_reset),
    .io_a(x369_sum_1_io_a),
    .io_b(x369_sum_1_io_b),
    .io_flow(x369_sum_1_io_flow),
    .io_result(x369_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@28450.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_57 ( // @[package.scala 93:22:@28462.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x255_sum x374_sum_1 ( // @[Math.scala 150:24:@28491.4]
    .clock(x374_sum_1_clock),
    .reset(x374_sum_1_reset),
    .io_a(x374_sum_1_io_a),
    .io_b(x374_sum_1_io_b),
    .io_flow(x374_sum_1_io_flow),
    .io_result(x374_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@28501.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_59 ( // @[package.scala 93:22:@28513.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  x377 x377_1 ( // @[Math.scala 262:24:@28536.4]
    .clock(x377_1_clock),
    .io_a(x377_1_io_a),
    .io_b(x377_1_io_b),
    .io_flow(x377_1_io_flow),
    .io_result(x377_1_io_result)
  );
  x377 x378_1 ( // @[Math.scala 262:24:@28548.4]
    .clock(x378_1_clock),
    .io_a(x378_1_io_a),
    .io_b(x378_1_io_b),
    .io_flow(x378_1_io_flow),
    .io_result(x378_1_io_result)
  );
  x377 x379_1 ( // @[Math.scala 262:24:@28560.4]
    .clock(x379_1_clock),
    .io_a(x379_1_io_a),
    .io_b(x379_1_io_b),
    .io_flow(x379_1_io_flow),
    .io_result(x379_1_io_result)
  );
  x377 x380_1 ( // @[Math.scala 262:24:@28572.4]
    .clock(x380_1_clock),
    .io_a(x380_1_io_a),
    .io_b(x380_1_io_b),
    .io_flow(x380_1_io_flow),
    .io_result(x380_1_io_result)
  );
  x377 x381_1 ( // @[Math.scala 262:24:@28584.4]
    .clock(x381_1_clock),
    .io_a(x381_1_io_a),
    .io_b(x381_1_io_b),
    .io_flow(x381_1_io_flow),
    .io_result(x381_1_io_result)
  );
  x377 x382_1 ( // @[Math.scala 262:24:@28596.4]
    .clock(x382_1_clock),
    .io_a(x382_1_io_a),
    .io_b(x382_1_io_b),
    .io_flow(x382_1_io_flow),
    .io_result(x382_1_io_result)
  );
  x377 x383_1 ( // @[Math.scala 262:24:@28608.4]
    .clock(x383_1_clock),
    .io_a(x383_1_io_a),
    .io_b(x383_1_io_b),
    .io_flow(x383_1_io_flow),
    .io_result(x383_1_io_result)
  );
  x377 x384_1 ( // @[Math.scala 262:24:@28620.4]
    .clock(x384_1_clock),
    .io_a(x384_1_io_a),
    .io_b(x384_1_io_b),
    .io_flow(x384_1_io_flow),
    .io_result(x384_1_io_result)
  );
  x377 x385_1 ( // @[Math.scala 262:24:@28632.4]
    .clock(x385_1_clock),
    .io_a(x385_1_io_a),
    .io_b(x385_1_io_b),
    .io_flow(x385_1_io_flow),
    .io_result(x385_1_io_result)
  );
  x386_x13 x386_x13_1 ( // @[Math.scala 150:24:@28642.4]
    .clock(x386_x13_1_clock),
    .reset(x386_x13_1_reset),
    .io_a(x386_x13_1_io_a),
    .io_b(x386_x13_1_io_b),
    .io_flow(x386_x13_1_io_flow),
    .io_result(x386_x13_1_io_result)
  );
  x386_x13 x387_x14_1 ( // @[Math.scala 150:24:@28652.4]
    .clock(x387_x14_1_clock),
    .reset(x387_x14_1_reset),
    .io_a(x387_x14_1_io_a),
    .io_b(x387_x14_1_io_b),
    .io_flow(x387_x14_1_io_flow),
    .io_result(x387_x14_1_io_result)
  );
  x386_x13 x388_x13_1 ( // @[Math.scala 150:24:@28662.4]
    .clock(x388_x13_1_clock),
    .reset(x388_x13_1_reset),
    .io_a(x388_x13_1_io_a),
    .io_b(x388_x13_1_io_b),
    .io_flow(x388_x13_1_io_flow),
    .io_result(x388_x13_1_io_result)
  );
  x386_x13 x389_x14_1 ( // @[Math.scala 150:24:@28672.4]
    .clock(x389_x14_1_clock),
    .reset(x389_x14_1_reset),
    .io_a(x389_x14_1_io_a),
    .io_b(x389_x14_1_io_b),
    .io_flow(x389_x14_1_io_flow),
    .io_result(x389_x14_1_io_result)
  );
  x386_x13 x390_x13_1 ( // @[Math.scala 150:24:@28682.4]
    .clock(x390_x13_1_clock),
    .reset(x390_x13_1_reset),
    .io_a(x390_x13_1_io_a),
    .io_b(x390_x13_1_io_b),
    .io_flow(x390_x13_1_io_flow),
    .io_result(x390_x13_1_io_result)
  );
  x386_x13 x391_x14_1 ( // @[Math.scala 150:24:@28692.4]
    .clock(x391_x14_1_clock),
    .reset(x391_x14_1_reset),
    .io_a(x391_x14_1_io_a),
    .io_b(x391_x14_1_io_b),
    .io_flow(x391_x14_1_io_flow),
    .io_result(x391_x14_1_io_result)
  );
  x386_x13 x392_x13_1 ( // @[Math.scala 150:24:@28702.4]
    .clock(x392_x13_1_clock),
    .reset(x392_x13_1_reset),
    .io_a(x392_x13_1_io_a),
    .io_b(x392_x13_1_io_b),
    .io_flow(x392_x13_1_io_flow),
    .io_result(x392_x13_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_60 ( // @[package.scala 93:22:@28712.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x386_x13 x393_sum_1 ( // @[Math.scala 150:24:@28721.4]
    .clock(x393_sum_1_clock),
    .reset(x393_sum_1_reset),
    .io_a(x393_sum_1_io_a),
    .io_b(x393_sum_1_io_b),
    .io_flow(x393_sum_1_io_flow),
    .io_result(x393_sum_1_io_result)
  );
  x394 x394_1 ( // @[Math.scala 720:24:@28731.4]
    .io_b(x394_1_io_b),
    .io_result(x394_1_io_result)
  );
  x395_mul x395_mul_1 ( // @[Math.scala 262:24:@28742.4]
    .clock(x395_mul_1_clock),
    .io_a(x395_mul_1_io_a),
    .io_b(x395_mul_1_io_b),
    .io_flow(x395_mul_1_io_flow),
    .io_result(x395_mul_1_io_result)
  );
  x396 x396_1 ( // @[Math.scala 720:24:@28752.4]
    .io_b(x396_1_io_b),
    .io_result(x396_1_io_result)
  );
  RetimeWrapper_253 RetimeWrapper_61 ( // @[package.scala 93:22:@28761.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x397_sub x397_sub_1 ( // @[Math.scala 191:24:@28770.4]
    .clock(x397_sub_1_clock),
    .reset(x397_sub_1_reset),
    .io_a(x397_sub_1_io_a),
    .io_b(x397_sub_1_io_b),
    .io_flow(x397_sub_1_io_flow),
    .io_result(x397_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@28783.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x397_sub x399_sub_1 ( // @[Math.scala 191:24:@28792.4]
    .clock(x399_sub_1_clock),
    .reset(x399_sub_1_reset),
    .io_a(x399_sub_1_io_a),
    .io_b(x399_sub_1_io_b),
    .io_flow(x399_sub_1_io_flow),
    .io_result(x399_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_63 ( // @[package.scala 93:22:@28805.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_64 ( // @[package.scala 93:22:@28817.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  x394 x403_1 ( // @[Math.scala 720:24:@28831.4]
    .io_b(x403_1_io_b),
    .io_result(x403_1_io_result)
  );
  x395_mul x404_mul_1 ( // @[Math.scala 262:24:@28842.4]
    .clock(x404_mul_1_clock),
    .io_a(x404_mul_1_io_a),
    .io_b(x404_mul_1_io_b),
    .io_flow(x404_mul_1_io_flow),
    .io_result(x404_mul_1_io_result)
  );
  x396 x405_1 ( // @[Math.scala 720:24:@28852.4]
    .io_b(x405_1_io_b),
    .io_result(x405_1_io_result)
  );
  RetimeWrapper_259 RetimeWrapper_65 ( // @[package.scala 93:22:@28861.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x386_x13 x406_sum_1 ( // @[Math.scala 150:24:@28870.4]
    .clock(x406_sum_1_clock),
    .reset(x406_sum_1_reset),
    .io_a(x406_sum_1_io_a),
    .io_b(x406_sum_1_io_b),
    .io_flow(x406_sum_1_io_flow),
    .io_result(x406_sum_1_io_result)
  );
  x377 x407_1 ( // @[Math.scala 262:24:@28882.4]
    .clock(x407_1_clock),
    .io_a(x407_1_io_a),
    .io_b(x407_1_io_b),
    .io_flow(x407_1_io_flow),
    .io_result(x407_1_io_result)
  );
  x377 x408_1 ( // @[Math.scala 262:24:@28894.4]
    .clock(x408_1_clock),
    .io_a(x408_1_io_a),
    .io_b(x408_1_io_b),
    .io_flow(x408_1_io_flow),
    .io_result(x408_1_io_result)
  );
  x377 x409_1 ( // @[Math.scala 262:24:@28906.4]
    .clock(x409_1_clock),
    .io_a(x409_1_io_a),
    .io_b(x409_1_io_b),
    .io_flow(x409_1_io_flow),
    .io_result(x409_1_io_result)
  );
  x377 x410_1 ( // @[Math.scala 262:24:@28918.4]
    .clock(x410_1_clock),
    .io_a(x410_1_io_a),
    .io_b(x410_1_io_b),
    .io_flow(x410_1_io_flow),
    .io_result(x410_1_io_result)
  );
  x377 x411_1 ( // @[Math.scala 262:24:@28930.4]
    .clock(x411_1_clock),
    .io_a(x411_1_io_a),
    .io_b(x411_1_io_b),
    .io_flow(x411_1_io_flow),
    .io_result(x411_1_io_result)
  );
  x377 x412_1 ( // @[Math.scala 262:24:@28942.4]
    .clock(x412_1_clock),
    .io_a(x412_1_io_a),
    .io_b(x412_1_io_b),
    .io_flow(x412_1_io_flow),
    .io_result(x412_1_io_result)
  );
  x377 x413_1 ( // @[Math.scala 262:24:@28954.4]
    .clock(x413_1_clock),
    .io_a(x413_1_io_a),
    .io_b(x413_1_io_b),
    .io_flow(x413_1_io_flow),
    .io_result(x413_1_io_result)
  );
  x377 x414_1 ( // @[Math.scala 262:24:@28966.4]
    .clock(x414_1_clock),
    .io_a(x414_1_io_a),
    .io_b(x414_1_io_b),
    .io_flow(x414_1_io_flow),
    .io_result(x414_1_io_result)
  );
  x377 x415_1 ( // @[Math.scala 262:24:@28978.4]
    .clock(x415_1_clock),
    .io_a(x415_1_io_a),
    .io_b(x415_1_io_b),
    .io_flow(x415_1_io_flow),
    .io_result(x415_1_io_result)
  );
  x386_x13 x416_x13_1 ( // @[Math.scala 150:24:@28990.4]
    .clock(x416_x13_1_clock),
    .reset(x416_x13_1_reset),
    .io_a(x416_x13_1_io_a),
    .io_b(x416_x13_1_io_b),
    .io_flow(x416_x13_1_io_flow),
    .io_result(x416_x13_1_io_result)
  );
  x386_x13 x417_x14_1 ( // @[Math.scala 150:24:@29000.4]
    .clock(x417_x14_1_clock),
    .reset(x417_x14_1_reset),
    .io_a(x417_x14_1_io_a),
    .io_b(x417_x14_1_io_b),
    .io_flow(x417_x14_1_io_flow),
    .io_result(x417_x14_1_io_result)
  );
  x386_x13 x418_x13_1 ( // @[Math.scala 150:24:@29010.4]
    .clock(x418_x13_1_clock),
    .reset(x418_x13_1_reset),
    .io_a(x418_x13_1_io_a),
    .io_b(x418_x13_1_io_b),
    .io_flow(x418_x13_1_io_flow),
    .io_result(x418_x13_1_io_result)
  );
  x386_x13 x419_x14_1 ( // @[Math.scala 150:24:@29020.4]
    .clock(x419_x14_1_clock),
    .reset(x419_x14_1_reset),
    .io_a(x419_x14_1_io_a),
    .io_b(x419_x14_1_io_b),
    .io_flow(x419_x14_1_io_flow),
    .io_result(x419_x14_1_io_result)
  );
  x386_x13 x420_x13_1 ( // @[Math.scala 150:24:@29030.4]
    .clock(x420_x13_1_clock),
    .reset(x420_x13_1_reset),
    .io_a(x420_x13_1_io_a),
    .io_b(x420_x13_1_io_b),
    .io_flow(x420_x13_1_io_flow),
    .io_result(x420_x13_1_io_result)
  );
  x386_x13 x421_x14_1 ( // @[Math.scala 150:24:@29040.4]
    .clock(x421_x14_1_clock),
    .reset(x421_x14_1_reset),
    .io_a(x421_x14_1_io_a),
    .io_b(x421_x14_1_io_b),
    .io_flow(x421_x14_1_io_flow),
    .io_result(x421_x14_1_io_result)
  );
  x386_x13 x422_x13_1 ( // @[Math.scala 150:24:@29050.4]
    .clock(x422_x13_1_clock),
    .reset(x422_x13_1_reset),
    .io_a(x422_x13_1_io_a),
    .io_b(x422_x13_1_io_b),
    .io_flow(x422_x13_1_io_flow),
    .io_result(x422_x13_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_66 ( // @[package.scala 93:22:@29060.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x386_x13 x423_sum_1 ( // @[Math.scala 150:24:@29069.4]
    .clock(x423_sum_1_clock),
    .reset(x423_sum_1_reset),
    .io_a(x423_sum_1_io_a),
    .io_b(x423_sum_1_io_b),
    .io_flow(x423_sum_1_io_flow),
    .io_result(x423_sum_1_io_result)
  );
  x394 x424_1 ( // @[Math.scala 720:24:@29079.4]
    .io_b(x424_1_io_b),
    .io_result(x424_1_io_result)
  );
  x395_mul x425_mul_1 ( // @[Math.scala 262:24:@29090.4]
    .clock(x425_mul_1_clock),
    .io_a(x425_mul_1_io_a),
    .io_b(x425_mul_1_io_b),
    .io_flow(x425_mul_1_io_flow),
    .io_result(x425_mul_1_io_result)
  );
  x396 x426_1 ( // @[Math.scala 720:24:@29100.4]
    .io_b(x426_1_io_b),
    .io_result(x426_1_io_result)
  );
  RetimeWrapper_253 RetimeWrapper_67 ( // @[package.scala 93:22:@29109.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x397_sub x427_sub_1 ( // @[Math.scala 191:24:@29118.4]
    .clock(x427_sub_1_clock),
    .reset(x427_sub_1_reset),
    .io_a(x427_sub_1_io_a),
    .io_b(x427_sub_1_io_b),
    .io_flow(x427_sub_1_io_flow),
    .io_result(x427_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_68 ( // @[package.scala 93:22:@29131.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  x397_sub x429_sub_1 ( // @[Math.scala 191:24:@29140.4]
    .clock(x429_sub_1_clock),
    .reset(x429_sub_1_reset),
    .io_a(x429_sub_1_io_a),
    .io_b(x429_sub_1_io_b),
    .io_flow(x429_sub_1_io_flow),
    .io_result(x429_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_69 ( // @[package.scala 93:22:@29153.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_70 ( // @[package.scala 93:22:@29165.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  x394 x433_1 ( // @[Math.scala 720:24:@29179.4]
    .io_b(x433_1_io_b),
    .io_result(x433_1_io_result)
  );
  x395_mul x434_mul_1 ( // @[Math.scala 262:24:@29190.4]
    .clock(x434_mul_1_clock),
    .io_a(x434_mul_1_io_a),
    .io_b(x434_mul_1_io_b),
    .io_flow(x434_mul_1_io_flow),
    .io_result(x434_mul_1_io_result)
  );
  x396 x435_1 ( // @[Math.scala 720:24:@29200.4]
    .io_b(x435_1_io_b),
    .io_result(x435_1_io_result)
  );
  RetimeWrapper_259 RetimeWrapper_71 ( // @[package.scala 93:22:@29209.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x386_x13 x436_sum_1 ( // @[Math.scala 150:24:@29218.4]
    .clock(x436_sum_1_clock),
    .reset(x436_sum_1_reset),
    .io_a(x436_sum_1_io_a),
    .io_b(x436_sum_1_io_b),
    .io_flow(x436_sum_1_io_flow),
    .io_result(x436_sum_1_io_result)
  );
  RetimeWrapper_278 RetimeWrapper_72 ( // @[package.scala 93:22:@29234.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_73 ( // @[package.scala 93:22:@29243.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_74 ( // @[package.scala 93:22:@29252.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_75 ( // @[package.scala 93:22:@29261.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  assign b274 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 62:18:@27069.4]
  assign b275 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 63:18:@27070.4]
  assign _T_205 = b274 & b275; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 67:30:@27072.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 67:37:@27073.4]
  assign _T_210 = io_in_x241_TID == 8'h0; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 69:76:@27078.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 69:62:@27079.4]
  assign _T_213 = io_in_x241_TDEST == 8'h0; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 69:101:@27080.4]
  assign x523_x276_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@27089.4 package.scala 96:25:@27090.4]
  assign b272_number = __io_result; // @[Math.scala 723:22:@27054.4 Math.scala 724:14:@27055.4]
  assign _T_243 = $signed(b272_number); // @[Math.scala 406:49:@27198.4]
  assign _T_245 = $signed(_T_243) & $signed(32'sh3); // @[Math.scala 406:56:@27200.4]
  assign _T_246 = $signed(_T_245); // @[Math.scala 406:56:@27201.4]
  assign x499_number = $unsigned(_T_246); // @[implicits.scala 133:21:@27202.4]
  assign _T_256 = $signed(x499_number); // @[Math.scala 406:49:@27211.4]
  assign _T_258 = $signed(_T_256) & $signed(32'sh3); // @[Math.scala 406:56:@27213.4]
  assign _T_259 = $signed(_T_258); // @[Math.scala 406:56:@27214.4]
  assign b273_number = __1_io_result; // @[Math.scala 723:22:@27066.4 Math.scala 724:14:@27067.4]
  assign _T_268 = $signed(b273_number); // @[Math.scala 406:49:@27222.4]
  assign _T_270 = $signed(_T_268) & $signed(32'sh3); // @[Math.scala 406:56:@27224.4]
  assign _T_271 = $signed(_T_270); // @[Math.scala 406:56:@27225.4]
  assign _T_275 = x499_number[31]; // @[FixedPoint.scala 50:25:@27231.4]
  assign _T_279 = _T_275 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27233.4]
  assign _T_280 = x499_number[31:2]; // @[FixedPoint.scala 18:52:@27234.4]
  assign _T_286 = _T_280 == 30'h3fffffff; // @[Math.scala 451:55:@27236.4]
  assign _T_287 = x499_number[1:0]; // @[FixedPoint.scala 18:52:@27237.4]
  assign _T_293 = _T_287 != 2'h0; // @[Math.scala 451:110:@27239.4]
  assign _T_294 = _T_286 & _T_293; // @[Math.scala 451:94:@27240.4]
  assign _T_296 = {_T_279,_T_280}; // @[Cat.scala 30:58:@27242.4]
  assign x284_1_number = _T_294 ? 32'h0 : _T_296; // @[Math.scala 454:20:@27243.4]
  assign _GEN_0 = {{9'd0}, x284_1_number}; // @[Math.scala 461:32:@27248.4]
  assign _T_301 = _GEN_0 << 9; // @[Math.scala 461:32:@27248.4]
  assign _GEN_1 = {{5'd0}, x284_1_number}; // @[Math.scala 461:32:@27253.4]
  assign _T_304 = _GEN_1 << 5; // @[Math.scala 461:32:@27253.4]
  assign _T_310 = b273_number[31]; // @[FixedPoint.scala 50:25:@27268.4]
  assign _T_314 = _T_310 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27270.4]
  assign _T_315 = b273_number[31:2]; // @[FixedPoint.scala 18:52:@27271.4]
  assign _T_321 = _T_315 == 30'h3fffffff; // @[Math.scala 451:55:@27273.4]
  assign _T_322 = b273_number[1:0]; // @[FixedPoint.scala 18:52:@27274.4]
  assign _T_328 = _T_322 != 2'h0; // @[Math.scala 451:110:@27276.4]
  assign _T_329 = _T_321 & _T_328; // @[Math.scala 451:94:@27277.4]
  assign _T_331 = {_T_314,_T_315}; // @[Cat.scala 30:58:@27279.4]
  assign _T_359 = ~ io_sigsIn_break; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:101:@27356.4]
  assign _T_363 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@27364.4 package.scala 96:25:@27365.4]
  assign _T_365 = io_rr ? _T_363 : 1'h0; // @[implicits.scala 55:10:@27366.4]
  assign _T_366 = _T_359 & _T_365; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:118:@27367.4]
  assign _T_368 = _T_366 & _T_359; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:206:@27369.4]
  assign _T_369 = _T_368 & io_sigsIn_backpressure; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:225:@27370.4]
  assign x528_b274_D3 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@27335.4 package.scala 96:25:@27336.4]
  assign _T_370 = _T_369 & x528_b274_D3; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 117:251:@27371.4]
  assign x526_b275_D3 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@27317.4 package.scala 96:25:@27318.4]
  assign x289_rdcol_number = x289_rdcol_1_io_result; // @[Math.scala 154:22:@27388.4 Math.scala 155:14:@27389.4]
  assign _T_387 = $signed(x289_rdcol_number); // @[Math.scala 406:49:@27397.4]
  assign _T_389 = $signed(_T_387) & $signed(32'sh3); // @[Math.scala 406:56:@27399.4]
  assign _T_390 = $signed(_T_389); // @[Math.scala 406:56:@27400.4]
  assign _T_394 = x289_rdcol_number[31]; // @[FixedPoint.scala 50:25:@27406.4]
  assign _T_398 = _T_394 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27408.4]
  assign _T_399 = x289_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@27409.4]
  assign _T_405 = _T_399 == 30'h3fffffff; // @[Math.scala 451:55:@27411.4]
  assign _T_406 = x289_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@27412.4]
  assign _T_412 = _T_406 != 2'h0; // @[Math.scala 451:110:@27414.4]
  assign _T_413 = _T_405 & _T_412; // @[Math.scala 451:94:@27415.4]
  assign _T_415 = {_T_398,_T_399}; // @[Cat.scala 30:58:@27417.4]
  assign _T_435 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@27466.4 package.scala 96:25:@27467.4]
  assign _T_437 = io_rr ? _T_435 : 1'h0; // @[implicits.scala 55:10:@27468.4]
  assign _T_438 = _T_359 & _T_437; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:118:@27469.4]
  assign _T_440 = _T_438 & _T_359; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:206:@27471.4]
  assign _T_441 = _T_440 & io_sigsIn_backpressure; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:225:@27472.4]
  assign _T_442 = _T_441 & x528_b274_D3; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 138:251:@27473.4]
  assign x534_b272_D6_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@27487.4 package.scala 96:25:@27488.4]
  assign _T_452 = $signed(x534_b272_D6_number); // @[Math.scala 476:37:@27493.4]
  assign x296 = $signed(_T_452) < $signed(32'sh0); // @[Math.scala 476:44:@27495.4]
  assign x535_x289_rdcol_D6_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@27503.4 package.scala 96:25:@27504.4]
  assign _T_463 = $signed(x535_x289_rdcol_D6_number); // @[Math.scala 476:37:@27509.4]
  assign x297 = $signed(_T_463) < $signed(32'sh0); // @[Math.scala 476:44:@27511.4]
  assign x536_x296_D1 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@27519.4 package.scala 96:25:@27520.4]
  assign x298 = x536_x296_D1 | x297; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 151:24:@27523.4]
  assign _T_502 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@27591.4 package.scala 96:25:@27592.4]
  assign _T_504 = io_rr ? _T_502 : 1'h0; // @[implicits.scala 55:10:@27593.4]
  assign _T_505 = _T_359 & _T_504; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 170:146:@27594.4]
  assign x541_x299_D2 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@27570.4 package.scala 96:25:@27571.4]
  assign _T_506 = _T_505 & x541_x299_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 170:234:@27595.4]
  assign x540_b274_D9 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@27561.4 package.scala 96:25:@27562.4]
  assign _T_507 = _T_506 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 170:242:@27596.4]
  assign x539_b275_D9 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@27552.4 package.scala 96:25:@27553.4]
  assign x543_b273_D6_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@27612.4 package.scala 96:25:@27613.4]
  assign _T_520 = $signed(x543_b273_D6_number); // @[Math.scala 476:37:@27620.4]
  assign x302 = $signed(_T_520) < $signed(32'sh0); // @[Math.scala 476:44:@27622.4]
  assign x303 = x296 | x302; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 186:59:@27625.4]
  assign _T_547 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@27666.4 package.scala 96:25:@27667.4]
  assign _T_549 = io_rr ? _T_547 : 1'h0; // @[implicits.scala 55:10:@27668.4]
  assign _T_550 = _T_359 & _T_549; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 199:194:@27669.4]
  assign x544_x304_D3 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@27636.4 package.scala 96:25:@27637.4]
  assign _T_551 = _T_550 & x544_x304_D3; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 199:282:@27670.4]
  assign _T_552 = _T_551 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 199:290:@27671.4]
  assign x307_rdcol_number = x307_rdcol_1_io_result; // @[Math.scala 154:22:@27690.4 Math.scala 155:14:@27691.4]
  assign _T_567 = $signed(x307_rdcol_number); // @[Math.scala 476:37:@27696.4]
  assign x308 = $signed(_T_567) < $signed(32'sh0); // @[Math.scala 476:44:@27698.4]
  assign x309 = x536_x296_D1 | x308; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 207:59:@27701.4]
  assign _T_583 = $signed(_T_567) & $signed(32'sh3); // @[Math.scala 406:56:@27712.4]
  assign _T_584 = $signed(_T_583); // @[Math.scala 406:56:@27713.4]
  assign _T_588 = x307_rdcol_number[31]; // @[FixedPoint.scala 50:25:@27719.4]
  assign _T_592 = _T_588 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27721.4]
  assign _T_593 = x307_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@27722.4]
  assign _T_599 = _T_593 == 30'h3fffffff; // @[Math.scala 451:55:@27724.4]
  assign _T_600 = x307_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@27725.4]
  assign _T_606 = _T_600 != 2'h0; // @[Math.scala 451:110:@27727.4]
  assign _T_607 = _T_599 & _T_606; // @[Math.scala 451:94:@27728.4]
  assign _T_609 = {_T_592,_T_593}; // @[Cat.scala 30:58:@27730.4]
  assign _T_638 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@27789.4 package.scala 96:25:@27790.4]
  assign _T_640 = io_rr ? _T_638 : 1'h0; // @[implicits.scala 55:10:@27791.4]
  assign _T_641 = _T_359 & _T_640; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 228:194:@27792.4]
  assign x549_x310_D2 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@27768.4 package.scala 96:25:@27769.4]
  assign _T_642 = _T_641 & x549_x310_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 228:282:@27793.4]
  assign _T_643 = _T_642 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 228:290:@27794.4]
  assign x316_rdcol_number = x316_rdcol_1_io_result; // @[Math.scala 154:22:@27813.4 Math.scala 155:14:@27814.4]
  assign _T_658 = $signed(x316_rdcol_number); // @[Math.scala 476:37:@27819.4]
  assign x317 = $signed(_T_658) < $signed(32'sh0); // @[Math.scala 476:44:@27821.4]
  assign x318 = x536_x296_D1 | x317; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 236:59:@27824.4]
  assign _T_674 = $signed(_T_658) & $signed(32'sh3); // @[Math.scala 406:56:@27835.4]
  assign _T_675 = $signed(_T_674); // @[Math.scala 406:56:@27836.4]
  assign _T_679 = x316_rdcol_number[31]; // @[FixedPoint.scala 50:25:@27842.4]
  assign _T_683 = _T_679 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27844.4]
  assign _T_684 = x316_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@27845.4]
  assign _T_690 = _T_684 == 30'h3fffffff; // @[Math.scala 451:55:@27847.4]
  assign _T_691 = x316_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@27848.4]
  assign _T_697 = _T_691 != 2'h0; // @[Math.scala 451:110:@27850.4]
  assign _T_698 = _T_690 & _T_697; // @[Math.scala 451:94:@27851.4]
  assign _T_700 = {_T_683,_T_684}; // @[Cat.scala 30:58:@27853.4]
  assign _T_726 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@27903.4 package.scala 96:25:@27904.4]
  assign _T_728 = io_rr ? _T_726 : 1'h0; // @[implicits.scala 55:10:@27905.4]
  assign _T_729 = _T_359 & _T_728; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 255:194:@27906.4]
  assign x552_x319_D2 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@27882.4 package.scala 96:25:@27883.4]
  assign _T_730 = _T_729 & x552_x319_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 255:282:@27907.4]
  assign _T_731 = _T_730 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 255:290:@27908.4]
  assign x325_rdrow_number = x325_rdrow_1_io_result; // @[Math.scala 195:22:@27927.4 Math.scala 196:14:@27928.4]
  assign _T_748 = $signed(x325_rdrow_number); // @[Math.scala 406:49:@27934.4]
  assign _T_750 = $signed(_T_748) & $signed(32'sh3); // @[Math.scala 406:56:@27936.4]
  assign _T_751 = $signed(_T_750); // @[Math.scala 406:56:@27937.4]
  assign x508_number = $unsigned(_T_751); // @[implicits.scala 133:21:@27938.4]
  assign x327 = $signed(_T_748) < $signed(32'sh0); // @[Math.scala 476:44:@27946.4]
  assign x328 = x327 | x297; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 265:24:@27949.4]
  assign _T_772 = $signed(x508_number); // @[Math.scala 406:49:@27958.4]
  assign _T_774 = $signed(_T_772) & $signed(32'sh3); // @[Math.scala 406:56:@27960.4]
  assign _T_775 = $signed(_T_774); // @[Math.scala 406:56:@27961.4]
  assign _T_779 = x508_number[31]; // @[FixedPoint.scala 50:25:@27967.4]
  assign _T_783 = _T_779 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27969.4]
  assign _T_784 = x508_number[31:2]; // @[FixedPoint.scala 18:52:@27970.4]
  assign _T_790 = _T_784 == 30'h3fffffff; // @[Math.scala 451:55:@27972.4]
  assign _T_791 = x508_number[1:0]; // @[FixedPoint.scala 18:52:@27973.4]
  assign _T_797 = _T_791 != 2'h0; // @[Math.scala 451:110:@27975.4]
  assign _T_798 = _T_790 & _T_797; // @[Math.scala 451:94:@27976.4]
  assign _T_800 = {_T_783,_T_784}; // @[Cat.scala 30:58:@27978.4]
  assign x331_1_number = _T_798 ? 32'h0 : _T_800; // @[Math.scala 454:20:@27979.4]
  assign _GEN_2 = {{9'd0}, x331_1_number}; // @[Math.scala 461:32:@27984.4]
  assign _T_805 = _GEN_2 << 9; // @[Math.scala 461:32:@27984.4]
  assign _GEN_3 = {{5'd0}, x331_1_number}; // @[Math.scala 461:32:@27989.4]
  assign _T_808 = _GEN_3 << 5; // @[Math.scala 461:32:@27989.4]
  assign _T_835 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@28048.4 package.scala 96:25:@28049.4]
  assign _T_837 = io_rr ? _T_835 : 1'h0; // @[implicits.scala 55:10:@28050.4]
  assign _T_838 = _T_359 & _T_837; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 290:194:@28051.4]
  assign x555_x329_D2 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@28027.4 package.scala 96:25:@28028.4]
  assign _T_839 = _T_838 & x555_x329_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 290:282:@28052.4]
  assign _T_840 = _T_839 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 290:290:@28053.4]
  assign x557_x302_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@28069.4 package.scala 96:25:@28070.4]
  assign x336 = x327 | x557_x302_D1; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 302:59:@28073.4]
  assign _T_872 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@28117.4 package.scala 96:25:@28118.4]
  assign _T_874 = io_rr ? _T_872 : 1'h0; // @[implicits.scala 55:10:@28119.4]
  assign _T_875 = _T_359 & _T_874; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 317:194:@28120.4]
  assign x559_x337_D2 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@28105.4 package.scala 96:25:@28106.4]
  assign _T_876 = _T_875 & x559_x337_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 317:282:@28121.4]
  assign _T_877 = _T_876 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 317:290:@28122.4]
  assign x341 = x327 | x308; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 321:59:@28133.4]
  assign _T_904 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@28175.4 package.scala 96:25:@28176.4]
  assign _T_906 = io_rr ? _T_904 : 1'h0; // @[implicits.scala 55:10:@28177.4]
  assign _T_907 = _T_359 & _T_906; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 334:194:@28178.4]
  assign x561_x342_D2 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@28163.4 package.scala 96:25:@28164.4]
  assign _T_908 = _T_907 & x561_x342_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 334:282:@28179.4]
  assign _T_909 = _T_908 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 334:290:@28180.4]
  assign x346 = x327 | x317; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 338:59:@28191.4]
  assign _T_936 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@28233.4 package.scala 96:25:@28234.4]
  assign _T_938 = io_rr ? _T_936 : 1'h0; // @[implicits.scala 55:10:@28235.4]
  assign _T_939 = _T_359 & _T_938; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 351:194:@28236.4]
  assign x563_x347_D2 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@28221.4 package.scala 96:25:@28222.4]
  assign _T_940 = _T_939 & x563_x347_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 351:282:@28237.4]
  assign _T_941 = _T_940 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 351:290:@28238.4]
  assign x351_rdrow_number = x351_rdrow_1_io_result; // @[Math.scala 195:22:@28257.4 Math.scala 196:14:@28258.4]
  assign _T_958 = $signed(x351_rdrow_number); // @[Math.scala 406:49:@28264.4]
  assign _T_960 = $signed(_T_958) & $signed(32'sh3); // @[Math.scala 406:56:@28266.4]
  assign _T_961 = $signed(_T_960); // @[Math.scala 406:56:@28267.4]
  assign x513_number = $unsigned(_T_961); // @[implicits.scala 133:21:@28268.4]
  assign x353 = $signed(_T_958) < $signed(32'sh0); // @[Math.scala 476:44:@28276.4]
  assign x354 = x353 | x297; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 361:24:@28279.4]
  assign _T_982 = $signed(x513_number); // @[Math.scala 406:49:@28288.4]
  assign _T_984 = $signed(_T_982) & $signed(32'sh3); // @[Math.scala 406:56:@28290.4]
  assign _T_985 = $signed(_T_984); // @[Math.scala 406:56:@28291.4]
  assign _T_989 = x513_number[31]; // @[FixedPoint.scala 50:25:@28297.4]
  assign _T_993 = _T_989 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28299.4]
  assign _T_994 = x513_number[31:2]; // @[FixedPoint.scala 18:52:@28300.4]
  assign _T_1000 = _T_994 == 30'h3fffffff; // @[Math.scala 451:55:@28302.4]
  assign _T_1001 = x513_number[1:0]; // @[FixedPoint.scala 18:52:@28303.4]
  assign _T_1007 = _T_1001 != 2'h0; // @[Math.scala 451:110:@28305.4]
  assign _T_1008 = _T_1000 & _T_1007; // @[Math.scala 451:94:@28306.4]
  assign _T_1010 = {_T_993,_T_994}; // @[Cat.scala 30:58:@28308.4]
  assign x357_1_number = _T_1008 ? 32'h0 : _T_1010; // @[Math.scala 454:20:@28309.4]
  assign _GEN_4 = {{9'd0}, x357_1_number}; // @[Math.scala 461:32:@28314.4]
  assign _T_1015 = _GEN_4 << 9; // @[Math.scala 461:32:@28314.4]
  assign _GEN_5 = {{5'd0}, x357_1_number}; // @[Math.scala 461:32:@28319.4]
  assign _T_1018 = _GEN_5 << 5; // @[Math.scala 461:32:@28319.4]
  assign _T_1042 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@28369.4 package.scala 96:25:@28370.4]
  assign _T_1044 = io_rr ? _T_1042 : 1'h0; // @[implicits.scala 55:10:@28371.4]
  assign _T_1045 = _T_359 & _T_1044; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 384:194:@28372.4]
  assign x565_x355_D2 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@28357.4 package.scala 96:25:@28358.4]
  assign _T_1046 = _T_1045 & x565_x355_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 384:282:@28373.4]
  assign _T_1047 = _T_1046 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 384:290:@28374.4]
  assign x362 = x353 | x557_x302_D1; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 388:24:@28385.4]
  assign _T_1071 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@28418.4 package.scala 96:25:@28419.4]
  assign _T_1073 = io_rr ? _T_1071 : 1'h0; // @[implicits.scala 55:10:@28420.4]
  assign _T_1074 = _T_359 & _T_1073; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 399:194:@28421.4]
  assign x566_x363_D2 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@28406.4 package.scala 96:25:@28407.4]
  assign _T_1075 = _T_1074 & x566_x363_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 399:282:@28422.4]
  assign _T_1076 = _T_1075 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 399:290:@28423.4]
  assign x367 = x353 | x308; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 403:24:@28434.4]
  assign _T_1100 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@28467.4 package.scala 96:25:@28468.4]
  assign _T_1102 = io_rr ? _T_1100 : 1'h0; // @[implicits.scala 55:10:@28469.4]
  assign _T_1103 = _T_359 & _T_1102; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 414:194:@28470.4]
  assign x567_x368_D2 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@28455.4 package.scala 96:25:@28456.4]
  assign _T_1104 = _T_1103 & x567_x368_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 414:282:@28471.4]
  assign _T_1105 = _T_1104 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 414:290:@28472.4]
  assign x372 = x353 | x317; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 424:59:@28483.4]
  assign _T_1131 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@28518.4 package.scala 96:25:@28519.4]
  assign _T_1133 = io_rr ? _T_1131 : 1'h0; // @[implicits.scala 55:10:@28520.4]
  assign _T_1134 = _T_359 & _T_1133; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 437:194:@28521.4]
  assign x568_x373_D2 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@28506.4 package.scala 96:25:@28507.4]
  assign _T_1135 = _T_1134 & x568_x373_D2; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 437:282:@28522.4]
  assign _T_1136 = _T_1135 & x540_b274_D9; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 437:290:@28523.4]
  assign x397_sub_number = x397_sub_1_io_result; // @[Math.scala 195:22:@28776.4 Math.scala 196:14:@28777.4]
  assign x399_sub_number = x399_sub_1_io_result; // @[Math.scala 195:22:@28798.4 Math.scala 196:14:@28799.4]
  assign x398 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@28788.4 package.scala 96:25:@28789.4]
  assign x400 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@28810.4 package.scala 96:25:@28811.4]
  assign x401 = x398 | x400; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 493:24:@28814.4]
  assign x571_x397_sub_D1_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@28822.4 package.scala 96:25:@28823.4]
  assign x427_sub_number = x427_sub_1_io_result; // @[Math.scala 195:22:@29124.4 Math.scala 196:14:@29125.4]
  assign x429_sub_number = x429_sub_1_io_result; // @[Math.scala 195:22:@29146.4 Math.scala 196:14:@29147.4]
  assign x428 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@29136.4 package.scala 96:25:@29137.4]
  assign x430 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@29158.4 package.scala 96:25:@29159.4]
  assign x431 = x428 | x430; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 569:24:@29162.4]
  assign x575_x427_sub_D1_number = RetimeWrapper_70_io_out; // @[package.scala 96:25:@29170.4 package.scala 96:25:@29171.4]
  assign x406_sum_number = x406_sum_1_io_result; // @[Math.scala 154:22:@28876.4 Math.scala 155:14:@28877.4]
  assign x436_sum_number = x436_sum_1_io_result; // @[Math.scala 154:22:@29224.4 Math.scala 155:14:@29225.4]
  assign _T_1478 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@29266.4 package.scala 96:25:@29267.4]
  assign _T_1480 = io_rr ? _T_1478 : 1'h0; // @[implicits.scala 55:10:@29268.4]
  assign x577_b274_D39 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@29248.4 package.scala 96:25:@29249.4]
  assign _T_1481 = _T_1480 & x577_b274_D39; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 593:117:@29269.4]
  assign x578_b275_D39 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@29257.4 package.scala 96:25:@29258.4]
  assign _T_1482 = _T_1481 & x578_b275_D39; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 593:123:@29270.4]
  assign x525_x500_D3_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@27308.4 package.scala 96:25:@27309.4]
  assign x529_x287_sum_D1_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@27344.4 package.scala 96:25:@27345.4]
  assign x530_x501_D3_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@27353.4 package.scala 96:25:@27354.4]
  assign x531_x293_sum_D1_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@27437.4 package.scala 96:25:@27438.4]
  assign x532_x505_D2_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@27446.4 package.scala 96:25:@27447.4]
  assign x537_x500_D9_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@27534.4 package.scala 96:25:@27535.4]
  assign x538_x293_sum_D7_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@27543.4 package.scala 96:25:@27544.4]
  assign x542_x505_D8_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@27579.4 package.scala 96:25:@27580.4]
  assign x545_x287_sum_D7_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@27645.4 package.scala 96:25:@27646.4]
  assign x546_x501_D9_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@27654.4 package.scala 96:25:@27655.4]
  assign x548_x313_sum_D1_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@27759.4 package.scala 96:25:@27760.4]
  assign x550_x506_D2_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@27777.4 package.scala 96:25:@27778.4]
  assign x551_x507_D2_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@27873.4 package.scala 96:25:@27874.4]
  assign x553_x322_sum_D1_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@27891.4 package.scala 96:25:@27892.4]
  assign x333_sum_number = x333_sum_1_io_result; // @[Math.scala 154:22:@28018.4 Math.scala 155:14:@28019.4]
  assign x556_x509_D2_number = RetimeWrapper_39_io_out; // @[package.scala 96:25:@28036.4 package.scala 96:25:@28037.4]
  assign x338_sum_number = x338_sum_1_io_result; // @[Math.scala 154:22:@28096.4 Math.scala 155:14:@28097.4]
  assign x343_sum_number = x343_sum_1_io_result; // @[Math.scala 154:22:@28154.4 Math.scala 155:14:@28155.4]
  assign x348_sum_number = x348_sum_1_io_result; // @[Math.scala 154:22:@28212.4 Math.scala 155:14:@28213.4]
  assign x359_sum_number = x359_sum_1_io_result; // @[Math.scala 154:22:@28339.4 Math.scala 155:14:@28340.4]
  assign x564_x514_D2_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@28348.4 package.scala 96:25:@28349.4]
  assign x364_sum_number = x364_sum_1_io_result; // @[Math.scala 154:22:@28397.4 Math.scala 155:14:@28398.4]
  assign x369_sum_number = x369_sum_1_io_result; // @[Math.scala 154:22:@28446.4 Math.scala 155:14:@28447.4]
  assign x374_sum_number = x374_sum_1_io_result; // @[Math.scala 154:22:@28497.4 Math.scala 155:14:@28498.4]
  assign io_in_x241_TREADY = _T_211 & _T_213; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 67:22:@27074.4 sm_x441_inr_Foreach_SAMPLER_BOX.scala 69:22:@27082.4]
  assign io_in_x242_TVALID = _T_1482 & io_sigsIn_backpressure; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 593:22:@29272.4]
  assign io_in_x242_TDATA = {{192'd0}, RetimeWrapper_72_io_out}; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 594:24:@29273.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@27052.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@27064.4]
  assign RetimeWrapper_clock = clock; // @[:@27085.4]
  assign RetimeWrapper_reset = reset; // @[:@27086.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27088.4]
  assign RetimeWrapper_io_in = io_in_x241_TDATA[63:0]; // @[package.scala 94:16:@27087.4]
  assign x278_lb_0_clock = clock; // @[:@27095.4]
  assign x278_lb_0_reset = reset; // @[:@27096.4]
  assign x278_lb_0_io_rPort_11_banks_1 = x546_x501_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@27674.4]
  assign x278_lb_0_io_rPort_11_banks_0 = x537_x500_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@27673.4]
  assign x278_lb_0_io_rPort_11_ofs_0 = x545_x287_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@27675.4]
  assign x278_lb_0_io_rPort_11_en_0 = _T_552 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@27677.4]
  assign x278_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27676.4]
  assign x278_lb_0_io_rPort_10_banks_1 = x542_x505_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@27599.4]
  assign x278_lb_0_io_rPort_10_banks_0 = x537_x500_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@27598.4]
  assign x278_lb_0_io_rPort_10_ofs_0 = x538_x293_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@27600.4]
  assign x278_lb_0_io_rPort_10_en_0 = _T_507 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@27602.4]
  assign x278_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27601.4]
  assign x278_lb_0_io_rPort_9_banks_1 = x550_x506_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27797.4]
  assign x278_lb_0_io_rPort_9_banks_0 = x537_x500_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@27796.4]
  assign x278_lb_0_io_rPort_9_ofs_0 = x548_x313_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@27798.4]
  assign x278_lb_0_io_rPort_9_en_0 = _T_643 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@27800.4]
  assign x278_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27799.4]
  assign x278_lb_0_io_rPort_8_banks_1 = x550_x506_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28475.4]
  assign x278_lb_0_io_rPort_8_banks_0 = x564_x514_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28474.4]
  assign x278_lb_0_io_rPort_8_ofs_0 = x369_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28476.4]
  assign x278_lb_0_io_rPort_8_en_0 = _T_1105 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28478.4]
  assign x278_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28477.4]
  assign x278_lb_0_io_rPort_7_banks_1 = x551_x507_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27911.4]
  assign x278_lb_0_io_rPort_7_banks_0 = x537_x500_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@27910.4]
  assign x278_lb_0_io_rPort_7_ofs_0 = x553_x322_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@27912.4]
  assign x278_lb_0_io_rPort_7_en_0 = _T_731 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@27914.4]
  assign x278_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27913.4]
  assign x278_lb_0_io_rPort_6_banks_1 = x551_x507_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28526.4]
  assign x278_lb_0_io_rPort_6_banks_0 = x564_x514_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28525.4]
  assign x278_lb_0_io_rPort_6_ofs_0 = x374_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28527.4]
  assign x278_lb_0_io_rPort_6_en_0 = _T_1136 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28529.4]
  assign x278_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28528.4]
  assign x278_lb_0_io_rPort_5_banks_1 = x542_x505_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@28377.4]
  assign x278_lb_0_io_rPort_5_banks_0 = x564_x514_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28376.4]
  assign x278_lb_0_io_rPort_5_ofs_0 = x359_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28378.4]
  assign x278_lb_0_io_rPort_5_en_0 = _T_1047 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28380.4]
  assign x278_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28379.4]
  assign x278_lb_0_io_rPort_4_banks_1 = x546_x501_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@28125.4]
  assign x278_lb_0_io_rPort_4_banks_0 = x556_x509_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28124.4]
  assign x278_lb_0_io_rPort_4_ofs_0 = x338_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28126.4]
  assign x278_lb_0_io_rPort_4_en_0 = _T_877 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28128.4]
  assign x278_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28127.4]
  assign x278_lb_0_io_rPort_3_banks_1 = x551_x507_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28241.4]
  assign x278_lb_0_io_rPort_3_banks_0 = x556_x509_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28240.4]
  assign x278_lb_0_io_rPort_3_ofs_0 = x348_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28242.4]
  assign x278_lb_0_io_rPort_3_en_0 = _T_941 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28244.4]
  assign x278_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28243.4]
  assign x278_lb_0_io_rPort_2_banks_1 = x542_x505_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@28056.4]
  assign x278_lb_0_io_rPort_2_banks_0 = x556_x509_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28055.4]
  assign x278_lb_0_io_rPort_2_ofs_0 = x333_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28057.4]
  assign x278_lb_0_io_rPort_2_en_0 = _T_840 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28059.4]
  assign x278_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28058.4]
  assign x278_lb_0_io_rPort_1_banks_1 = x550_x506_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28183.4]
  assign x278_lb_0_io_rPort_1_banks_0 = x556_x509_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28182.4]
  assign x278_lb_0_io_rPort_1_ofs_0 = x343_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28184.4]
  assign x278_lb_0_io_rPort_1_en_0 = _T_909 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28186.4]
  assign x278_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28185.4]
  assign x278_lb_0_io_rPort_0_banks_1 = x546_x501_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@28426.4]
  assign x278_lb_0_io_rPort_0_banks_0 = x564_x514_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@28425.4]
  assign x278_lb_0_io_rPort_0_ofs_0 = x364_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@28427.4]
  assign x278_lb_0_io_rPort_0_en_0 = _T_1076 & x539_b275_D9; // @[MemInterfaceType.scala 110:79:@28429.4]
  assign x278_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28428.4]
  assign x278_lb_0_io_wPort_1_banks_1 = x532_x505_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@27476.4]
  assign x278_lb_0_io_wPort_1_banks_0 = x525_x500_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@27475.4]
  assign x278_lb_0_io_wPort_1_ofs_0 = x531_x293_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@27477.4]
  assign x278_lb_0_io_wPort_1_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@27478.4]
  assign x278_lb_0_io_wPort_1_en_0 = _T_442 & x526_b275_D3; // @[MemInterfaceType.scala 93:57:@27480.4]
  assign x278_lb_0_io_wPort_0_banks_1 = x530_x501_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@27374.4]
  assign x278_lb_0_io_wPort_0_banks_0 = x525_x500_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@27373.4]
  assign x278_lb_0_io_wPort_0_ofs_0 = x529_x287_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@27375.4]
  assign x278_lb_0_io_wPort_0_data_0 = RetimeWrapper_4_io_out; // @[MemInterfaceType.scala 90:56:@27376.4]
  assign x278_lb_0_io_wPort_0_en_0 = _T_370 & x526_b275_D3; // @[MemInterfaceType.scala 93:57:@27378.4]
  assign x504_sub_1_clock = clock; // @[:@27258.4]
  assign x504_sub_1_reset = reset; // @[:@27259.4]
  assign x504_sub_1_io_a = _T_301[31:0]; // @[Math.scala 192:17:@27260.4]
  assign x504_sub_1_io_b = _T_304[31:0]; // @[Math.scala 193:17:@27261.4]
  assign x504_sub_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@27262.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27285.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27286.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27288.4]
  assign RetimeWrapper_1_io_in = _T_329 ? 32'h0 : _T_331; // @[package.scala 94:16:@27287.4]
  assign x287_sum_1_clock = clock; // @[:@27294.4]
  assign x287_sum_1_reset = reset; // @[:@27295.4]
  assign x287_sum_1_io_a = x504_sub_1_io_result; // @[Math.scala 151:17:@27296.4]
  assign x287_sum_1_io_b = RetimeWrapper_1_io_out; // @[Math.scala 152:17:@27297.4]
  assign x287_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@27298.4]
  assign RetimeWrapper_2_clock = clock; // @[:@27304.4]
  assign RetimeWrapper_2_reset = reset; // @[:@27305.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27307.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_259); // @[package.scala 94:16:@27306.4]
  assign RetimeWrapper_3_clock = clock; // @[:@27313.4]
  assign RetimeWrapper_3_reset = reset; // @[:@27314.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27316.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27315.4]
  assign RetimeWrapper_4_clock = clock; // @[:@27322.4]
  assign RetimeWrapper_4_reset = reset; // @[:@27323.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27325.4]
  assign RetimeWrapper_4_io_in = x523_x276_D1_0_number[31:0]; // @[package.scala 94:16:@27324.4]
  assign RetimeWrapper_5_clock = clock; // @[:@27331.4]
  assign RetimeWrapper_5_reset = reset; // @[:@27332.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27334.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27333.4]
  assign RetimeWrapper_6_clock = clock; // @[:@27340.4]
  assign RetimeWrapper_6_reset = reset; // @[:@27341.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27343.4]
  assign RetimeWrapper_6_io_in = x287_sum_1_io_result; // @[package.scala 94:16:@27342.4]
  assign RetimeWrapper_7_clock = clock; // @[:@27349.4]
  assign RetimeWrapper_7_reset = reset; // @[:@27350.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27352.4]
  assign RetimeWrapper_7_io_in = $unsigned(_T_271); // @[package.scala 94:16:@27351.4]
  assign RetimeWrapper_8_clock = clock; // @[:@27360.4]
  assign RetimeWrapper_8_reset = reset; // @[:@27361.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27363.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27362.4]
  assign x289_rdcol_1_clock = clock; // @[:@27383.4]
  assign x289_rdcol_1_reset = reset; // @[:@27384.4]
  assign x289_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@27385.4]
  assign x289_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@27386.4]
  assign x289_rdcol_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@27387.4]
  assign x293_sum_1_clock = clock; // @[:@27423.4]
  assign x293_sum_1_reset = reset; // @[:@27424.4]
  assign x293_sum_1_io_a = x504_sub_1_io_result; // @[Math.scala 151:17:@27425.4]
  assign x293_sum_1_io_b = _T_413 ? 32'h0 : _T_415; // @[Math.scala 152:17:@27426.4]
  assign x293_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@27427.4]
  assign RetimeWrapper_9_clock = clock; // @[:@27433.4]
  assign RetimeWrapper_9_reset = reset; // @[:@27434.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27436.4]
  assign RetimeWrapper_9_io_in = x293_sum_1_io_result; // @[package.scala 94:16:@27435.4]
  assign RetimeWrapper_10_clock = clock; // @[:@27442.4]
  assign RetimeWrapper_10_reset = reset; // @[:@27443.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27445.4]
  assign RetimeWrapper_10_io_in = $unsigned(_T_390); // @[package.scala 94:16:@27444.4]
  assign RetimeWrapper_11_clock = clock; // @[:@27451.4]
  assign RetimeWrapper_11_reset = reset; // @[:@27452.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27454.4]
  assign RetimeWrapper_11_io_in = x523_x276_D1_0_number[63:32]; // @[package.scala 94:16:@27453.4]
  assign RetimeWrapper_12_clock = clock; // @[:@27462.4]
  assign RetimeWrapper_12_reset = reset; // @[:@27463.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27465.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27464.4]
  assign RetimeWrapper_13_clock = clock; // @[:@27483.4]
  assign RetimeWrapper_13_reset = reset; // @[:@27484.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27486.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@27485.4]
  assign RetimeWrapper_14_clock = clock; // @[:@27499.4]
  assign RetimeWrapper_14_reset = reset; // @[:@27500.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27502.4]
  assign RetimeWrapper_14_io_in = x289_rdcol_1_io_result; // @[package.scala 94:16:@27501.4]
  assign RetimeWrapper_15_clock = clock; // @[:@27515.4]
  assign RetimeWrapper_15_reset = reset; // @[:@27516.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27518.4]
  assign RetimeWrapper_15_io_in = $signed(_T_452) < $signed(32'sh0); // @[package.scala 94:16:@27517.4]
  assign RetimeWrapper_16_clock = clock; // @[:@27530.4]
  assign RetimeWrapper_16_reset = reset; // @[:@27531.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27533.4]
  assign RetimeWrapper_16_io_in = $unsigned(_T_259); // @[package.scala 94:16:@27532.4]
  assign RetimeWrapper_17_clock = clock; // @[:@27539.4]
  assign RetimeWrapper_17_reset = reset; // @[:@27540.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27542.4]
  assign RetimeWrapper_17_io_in = x293_sum_1_io_result; // @[package.scala 94:16:@27541.4]
  assign RetimeWrapper_18_clock = clock; // @[:@27548.4]
  assign RetimeWrapper_18_reset = reset; // @[:@27549.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27551.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27550.4]
  assign RetimeWrapper_19_clock = clock; // @[:@27557.4]
  assign RetimeWrapper_19_reset = reset; // @[:@27558.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27560.4]
  assign RetimeWrapper_19_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27559.4]
  assign RetimeWrapper_20_clock = clock; // @[:@27566.4]
  assign RetimeWrapper_20_reset = reset; // @[:@27567.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27569.4]
  assign RetimeWrapper_20_io_in = ~ x298; // @[package.scala 94:16:@27568.4]
  assign RetimeWrapper_21_clock = clock; // @[:@27575.4]
  assign RetimeWrapper_21_reset = reset; // @[:@27576.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27578.4]
  assign RetimeWrapper_21_io_in = $unsigned(_T_390); // @[package.scala 94:16:@27577.4]
  assign RetimeWrapper_22_clock = clock; // @[:@27587.4]
  assign RetimeWrapper_22_reset = reset; // @[:@27588.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27590.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27589.4]
  assign RetimeWrapper_23_clock = clock; // @[:@27608.4]
  assign RetimeWrapper_23_reset = reset; // @[:@27609.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27611.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@27610.4]
  assign RetimeWrapper_24_clock = clock; // @[:@27632.4]
  assign RetimeWrapper_24_reset = reset; // @[:@27633.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27635.4]
  assign RetimeWrapper_24_io_in = ~ x303; // @[package.scala 94:16:@27634.4]
  assign RetimeWrapper_25_clock = clock; // @[:@27641.4]
  assign RetimeWrapper_25_reset = reset; // @[:@27642.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27644.4]
  assign RetimeWrapper_25_io_in = x287_sum_1_io_result; // @[package.scala 94:16:@27643.4]
  assign RetimeWrapper_26_clock = clock; // @[:@27650.4]
  assign RetimeWrapper_26_reset = reset; // @[:@27651.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27653.4]
  assign RetimeWrapper_26_io_in = $unsigned(_T_271); // @[package.scala 94:16:@27652.4]
  assign RetimeWrapper_27_clock = clock; // @[:@27662.4]
  assign RetimeWrapper_27_reset = reset; // @[:@27663.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27665.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27664.4]
  assign x307_rdcol_1_clock = clock; // @[:@27685.4]
  assign x307_rdcol_1_reset = reset; // @[:@27686.4]
  assign x307_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@27687.4]
  assign x307_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@27688.4]
  assign x307_rdcol_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@27689.4]
  assign RetimeWrapper_28_clock = clock; // @[:@27736.4]
  assign RetimeWrapper_28_reset = reset; // @[:@27737.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27739.4]
  assign RetimeWrapper_28_io_in = x504_sub_1_io_result; // @[package.scala 94:16:@27738.4]
  assign x313_sum_1_clock = clock; // @[:@27745.4]
  assign x313_sum_1_reset = reset; // @[:@27746.4]
  assign x313_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@27747.4]
  assign x313_sum_1_io_b = _T_607 ? 32'h0 : _T_609; // @[Math.scala 152:17:@27748.4]
  assign x313_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@27749.4]
  assign RetimeWrapper_29_clock = clock; // @[:@27755.4]
  assign RetimeWrapper_29_reset = reset; // @[:@27756.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27758.4]
  assign RetimeWrapper_29_io_in = x313_sum_1_io_result; // @[package.scala 94:16:@27757.4]
  assign RetimeWrapper_30_clock = clock; // @[:@27764.4]
  assign RetimeWrapper_30_reset = reset; // @[:@27765.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27767.4]
  assign RetimeWrapper_30_io_in = ~ x309; // @[package.scala 94:16:@27766.4]
  assign RetimeWrapper_31_clock = clock; // @[:@27773.4]
  assign RetimeWrapper_31_reset = reset; // @[:@27774.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27776.4]
  assign RetimeWrapper_31_io_in = $unsigned(_T_584); // @[package.scala 94:16:@27775.4]
  assign RetimeWrapper_32_clock = clock; // @[:@27785.4]
  assign RetimeWrapper_32_reset = reset; // @[:@27786.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27788.4]
  assign RetimeWrapper_32_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27787.4]
  assign x316_rdcol_1_clock = clock; // @[:@27808.4]
  assign x316_rdcol_1_reset = reset; // @[:@27809.4]
  assign x316_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@27810.4]
  assign x316_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@27811.4]
  assign x316_rdcol_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@27812.4]
  assign x322_sum_1_clock = clock; // @[:@27859.4]
  assign x322_sum_1_reset = reset; // @[:@27860.4]
  assign x322_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@27861.4]
  assign x322_sum_1_io_b = _T_698 ? 32'h0 : _T_700; // @[Math.scala 152:17:@27862.4]
  assign x322_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@27863.4]
  assign RetimeWrapper_33_clock = clock; // @[:@27869.4]
  assign RetimeWrapper_33_reset = reset; // @[:@27870.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27872.4]
  assign RetimeWrapper_33_io_in = $unsigned(_T_675); // @[package.scala 94:16:@27871.4]
  assign RetimeWrapper_34_clock = clock; // @[:@27878.4]
  assign RetimeWrapper_34_reset = reset; // @[:@27879.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27881.4]
  assign RetimeWrapper_34_io_in = ~ x318; // @[package.scala 94:16:@27880.4]
  assign RetimeWrapper_35_clock = clock; // @[:@27887.4]
  assign RetimeWrapper_35_reset = reset; // @[:@27888.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27890.4]
  assign RetimeWrapper_35_io_in = x322_sum_1_io_result; // @[package.scala 94:16:@27889.4]
  assign RetimeWrapper_36_clock = clock; // @[:@27899.4]
  assign RetimeWrapper_36_reset = reset; // @[:@27900.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27902.4]
  assign RetimeWrapper_36_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27901.4]
  assign x325_rdrow_1_clock = clock; // @[:@27922.4]
  assign x325_rdrow_1_reset = reset; // @[:@27923.4]
  assign x325_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@27924.4]
  assign x325_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@27925.4]
  assign x325_rdrow_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@27926.4]
  assign x512_sub_1_clock = clock; // @[:@27994.4]
  assign x512_sub_1_reset = reset; // @[:@27995.4]
  assign x512_sub_1_io_a = _T_805[31:0]; // @[Math.scala 192:17:@27996.4]
  assign x512_sub_1_io_b = _T_808[31:0]; // @[Math.scala 193:17:@27997.4]
  assign x512_sub_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@27998.4]
  assign RetimeWrapper_37_clock = clock; // @[:@28004.4]
  assign RetimeWrapper_37_reset = reset; // @[:@28005.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28007.4]
  assign RetimeWrapper_37_io_in = _T_413 ? 32'h0 : _T_415; // @[package.scala 94:16:@28006.4]
  assign x333_sum_1_clock = clock; // @[:@28013.4]
  assign x333_sum_1_reset = reset; // @[:@28014.4]
  assign x333_sum_1_io_a = x512_sub_1_io_result; // @[Math.scala 151:17:@28015.4]
  assign x333_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@28016.4]
  assign x333_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28017.4]
  assign RetimeWrapper_38_clock = clock; // @[:@28023.4]
  assign RetimeWrapper_38_reset = reset; // @[:@28024.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28026.4]
  assign RetimeWrapper_38_io_in = ~ x328; // @[package.scala 94:16:@28025.4]
  assign RetimeWrapper_39_clock = clock; // @[:@28032.4]
  assign RetimeWrapper_39_reset = reset; // @[:@28033.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28035.4]
  assign RetimeWrapper_39_io_in = $unsigned(_T_775); // @[package.scala 94:16:@28034.4]
  assign RetimeWrapper_40_clock = clock; // @[:@28044.4]
  assign RetimeWrapper_40_reset = reset; // @[:@28045.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28047.4]
  assign RetimeWrapper_40_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28046.4]
  assign RetimeWrapper_41_clock = clock; // @[:@28065.4]
  assign RetimeWrapper_41_reset = reset; // @[:@28066.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28068.4]
  assign RetimeWrapper_41_io_in = $signed(_T_520) < $signed(32'sh0); // @[package.scala 94:16:@28067.4]
  assign RetimeWrapper_42_clock = clock; // @[:@28080.4]
  assign RetimeWrapper_42_reset = reset; // @[:@28081.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28083.4]
  assign RetimeWrapper_42_io_in = _T_329 ? 32'h0 : _T_331; // @[package.scala 94:16:@28082.4]
  assign x338_sum_1_clock = clock; // @[:@28091.4]
  assign x338_sum_1_reset = reset; // @[:@28092.4]
  assign x338_sum_1_io_a = x512_sub_1_io_result; // @[Math.scala 151:17:@28093.4]
  assign x338_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@28094.4]
  assign x338_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28095.4]
  assign RetimeWrapper_43_clock = clock; // @[:@28101.4]
  assign RetimeWrapper_43_reset = reset; // @[:@28102.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28104.4]
  assign RetimeWrapper_43_io_in = ~ x336; // @[package.scala 94:16:@28103.4]
  assign RetimeWrapper_44_clock = clock; // @[:@28113.4]
  assign RetimeWrapper_44_reset = reset; // @[:@28114.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28116.4]
  assign RetimeWrapper_44_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28115.4]
  assign RetimeWrapper_45_clock = clock; // @[:@28140.4]
  assign RetimeWrapper_45_reset = reset; // @[:@28141.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28143.4]
  assign RetimeWrapper_45_io_in = _T_607 ? 32'h0 : _T_609; // @[package.scala 94:16:@28142.4]
  assign x343_sum_1_clock = clock; // @[:@28149.4]
  assign x343_sum_1_reset = reset; // @[:@28150.4]
  assign x343_sum_1_io_a = x512_sub_1_io_result; // @[Math.scala 151:17:@28151.4]
  assign x343_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@28152.4]
  assign x343_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28153.4]
  assign RetimeWrapper_46_clock = clock; // @[:@28159.4]
  assign RetimeWrapper_46_reset = reset; // @[:@28160.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28162.4]
  assign RetimeWrapper_46_io_in = ~ x341; // @[package.scala 94:16:@28161.4]
  assign RetimeWrapper_47_clock = clock; // @[:@28171.4]
  assign RetimeWrapper_47_reset = reset; // @[:@28172.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28174.4]
  assign RetimeWrapper_47_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28173.4]
  assign RetimeWrapper_48_clock = clock; // @[:@28198.4]
  assign RetimeWrapper_48_reset = reset; // @[:@28199.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28201.4]
  assign RetimeWrapper_48_io_in = _T_698 ? 32'h0 : _T_700; // @[package.scala 94:16:@28200.4]
  assign x348_sum_1_clock = clock; // @[:@28207.4]
  assign x348_sum_1_reset = reset; // @[:@28208.4]
  assign x348_sum_1_io_a = x512_sub_1_io_result; // @[Math.scala 151:17:@28209.4]
  assign x348_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@28210.4]
  assign x348_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28211.4]
  assign RetimeWrapper_49_clock = clock; // @[:@28217.4]
  assign RetimeWrapper_49_reset = reset; // @[:@28218.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28220.4]
  assign RetimeWrapper_49_io_in = ~ x346; // @[package.scala 94:16:@28219.4]
  assign RetimeWrapper_50_clock = clock; // @[:@28229.4]
  assign RetimeWrapper_50_reset = reset; // @[:@28230.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28232.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28231.4]
  assign x351_rdrow_1_clock = clock; // @[:@28252.4]
  assign x351_rdrow_1_reset = reset; // @[:@28253.4]
  assign x351_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@28254.4]
  assign x351_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@28255.4]
  assign x351_rdrow_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@28256.4]
  assign x517_sub_1_clock = clock; // @[:@28324.4]
  assign x517_sub_1_reset = reset; // @[:@28325.4]
  assign x517_sub_1_io_a = _T_1015[31:0]; // @[Math.scala 192:17:@28326.4]
  assign x517_sub_1_io_b = _T_1018[31:0]; // @[Math.scala 193:17:@28327.4]
  assign x517_sub_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@28328.4]
  assign x359_sum_1_clock = clock; // @[:@28334.4]
  assign x359_sum_1_reset = reset; // @[:@28335.4]
  assign x359_sum_1_io_a = x517_sub_1_io_result; // @[Math.scala 151:17:@28336.4]
  assign x359_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@28337.4]
  assign x359_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28338.4]
  assign RetimeWrapper_51_clock = clock; // @[:@28344.4]
  assign RetimeWrapper_51_reset = reset; // @[:@28345.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28347.4]
  assign RetimeWrapper_51_io_in = $unsigned(_T_985); // @[package.scala 94:16:@28346.4]
  assign RetimeWrapper_52_clock = clock; // @[:@28353.4]
  assign RetimeWrapper_52_reset = reset; // @[:@28354.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28356.4]
  assign RetimeWrapper_52_io_in = ~ x354; // @[package.scala 94:16:@28355.4]
  assign RetimeWrapper_53_clock = clock; // @[:@28365.4]
  assign RetimeWrapper_53_reset = reset; // @[:@28366.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28368.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28367.4]
  assign x364_sum_1_clock = clock; // @[:@28392.4]
  assign x364_sum_1_reset = reset; // @[:@28393.4]
  assign x364_sum_1_io_a = x517_sub_1_io_result; // @[Math.scala 151:17:@28394.4]
  assign x364_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@28395.4]
  assign x364_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28396.4]
  assign RetimeWrapper_54_clock = clock; // @[:@28402.4]
  assign RetimeWrapper_54_reset = reset; // @[:@28403.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28405.4]
  assign RetimeWrapper_54_io_in = ~ x362; // @[package.scala 94:16:@28404.4]
  assign RetimeWrapper_55_clock = clock; // @[:@28414.4]
  assign RetimeWrapper_55_reset = reset; // @[:@28415.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28417.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28416.4]
  assign x369_sum_1_clock = clock; // @[:@28441.4]
  assign x369_sum_1_reset = reset; // @[:@28442.4]
  assign x369_sum_1_io_a = x517_sub_1_io_result; // @[Math.scala 151:17:@28443.4]
  assign x369_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@28444.4]
  assign x369_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28445.4]
  assign RetimeWrapper_56_clock = clock; // @[:@28451.4]
  assign RetimeWrapper_56_reset = reset; // @[:@28452.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28454.4]
  assign RetimeWrapper_56_io_in = ~ x367; // @[package.scala 94:16:@28453.4]
  assign RetimeWrapper_57_clock = clock; // @[:@28463.4]
  assign RetimeWrapper_57_reset = reset; // @[:@28464.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28466.4]
  assign RetimeWrapper_57_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28465.4]
  assign x374_sum_1_clock = clock; // @[:@28492.4]
  assign x374_sum_1_reset = reset; // @[:@28493.4]
  assign x374_sum_1_io_a = x517_sub_1_io_result; // @[Math.scala 151:17:@28494.4]
  assign x374_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@28495.4]
  assign x374_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28496.4]
  assign RetimeWrapper_58_clock = clock; // @[:@28502.4]
  assign RetimeWrapper_58_reset = reset; // @[:@28503.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28505.4]
  assign RetimeWrapper_58_io_in = ~ x372; // @[package.scala 94:16:@28504.4]
  assign RetimeWrapper_59_clock = clock; // @[:@28514.4]
  assign RetimeWrapper_59_reset = reset; // @[:@28515.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28517.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28516.4]
  assign x377_1_clock = clock; // @[:@28537.4]
  assign x377_1_io_a = x278_lb_0_io_rPort_10_output_0; // @[Math.scala 263:17:@28539.4]
  assign x377_1_io_b = 32'h1; // @[Math.scala 264:17:@28540.4]
  assign x377_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28541.4]
  assign x378_1_clock = clock; // @[:@28549.4]
  assign x378_1_io_a = x278_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@28551.4]
  assign x378_1_io_b = 32'h2; // @[Math.scala 264:17:@28552.4]
  assign x378_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28553.4]
  assign x379_1_clock = clock; // @[:@28561.4]
  assign x379_1_io_a = x278_lb_0_io_rPort_9_output_0; // @[Math.scala 263:17:@28563.4]
  assign x379_1_io_b = 32'h1; // @[Math.scala 264:17:@28564.4]
  assign x379_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28565.4]
  assign x380_1_clock = clock; // @[:@28573.4]
  assign x380_1_io_a = x278_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@28575.4]
  assign x380_1_io_b = 32'h2; // @[Math.scala 264:17:@28576.4]
  assign x380_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28577.4]
  assign x381_1_clock = clock; // @[:@28585.4]
  assign x381_1_io_a = x278_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@28587.4]
  assign x381_1_io_b = 32'h4; // @[Math.scala 264:17:@28588.4]
  assign x381_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28589.4]
  assign x382_1_clock = clock; // @[:@28597.4]
  assign x382_1_io_a = x278_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@28599.4]
  assign x382_1_io_b = 32'h2; // @[Math.scala 264:17:@28600.4]
  assign x382_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28601.4]
  assign x383_1_clock = clock; // @[:@28609.4]
  assign x383_1_io_a = x278_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@28611.4]
  assign x383_1_io_b = 32'h1; // @[Math.scala 264:17:@28612.4]
  assign x383_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28613.4]
  assign x384_1_clock = clock; // @[:@28621.4]
  assign x384_1_io_a = x278_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@28623.4]
  assign x384_1_io_b = 32'h2; // @[Math.scala 264:17:@28624.4]
  assign x384_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28625.4]
  assign x385_1_clock = clock; // @[:@28633.4]
  assign x385_1_io_a = x278_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@28635.4]
  assign x385_1_io_b = 32'h1; // @[Math.scala 264:17:@28636.4]
  assign x385_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28637.4]
  assign x386_x13_1_clock = clock; // @[:@28643.4]
  assign x386_x13_1_reset = reset; // @[:@28644.4]
  assign x386_x13_1_io_a = x377_1_io_result; // @[Math.scala 151:17:@28645.4]
  assign x386_x13_1_io_b = x378_1_io_result; // @[Math.scala 152:17:@28646.4]
  assign x386_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28647.4]
  assign x387_x14_1_clock = clock; // @[:@28653.4]
  assign x387_x14_1_reset = reset; // @[:@28654.4]
  assign x387_x14_1_io_a = x379_1_io_result; // @[Math.scala 151:17:@28655.4]
  assign x387_x14_1_io_b = x380_1_io_result; // @[Math.scala 152:17:@28656.4]
  assign x387_x14_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28657.4]
  assign x388_x13_1_clock = clock; // @[:@28663.4]
  assign x388_x13_1_reset = reset; // @[:@28664.4]
  assign x388_x13_1_io_a = x381_1_io_result; // @[Math.scala 151:17:@28665.4]
  assign x388_x13_1_io_b = x382_1_io_result; // @[Math.scala 152:17:@28666.4]
  assign x388_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28667.4]
  assign x389_x14_1_clock = clock; // @[:@28673.4]
  assign x389_x14_1_reset = reset; // @[:@28674.4]
  assign x389_x14_1_io_a = x383_1_io_result; // @[Math.scala 151:17:@28675.4]
  assign x389_x14_1_io_b = x384_1_io_result; // @[Math.scala 152:17:@28676.4]
  assign x389_x14_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28677.4]
  assign x390_x13_1_clock = clock; // @[:@28683.4]
  assign x390_x13_1_reset = reset; // @[:@28684.4]
  assign x390_x13_1_io_a = x386_x13_1_io_result; // @[Math.scala 151:17:@28685.4]
  assign x390_x13_1_io_b = x387_x14_1_io_result; // @[Math.scala 152:17:@28686.4]
  assign x390_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28687.4]
  assign x391_x14_1_clock = clock; // @[:@28693.4]
  assign x391_x14_1_reset = reset; // @[:@28694.4]
  assign x391_x14_1_io_a = x388_x13_1_io_result; // @[Math.scala 151:17:@28695.4]
  assign x391_x14_1_io_b = x389_x14_1_io_result; // @[Math.scala 152:17:@28696.4]
  assign x391_x14_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28697.4]
  assign x392_x13_1_clock = clock; // @[:@28703.4]
  assign x392_x13_1_reset = reset; // @[:@28704.4]
  assign x392_x13_1_io_a = x390_x13_1_io_result; // @[Math.scala 151:17:@28705.4]
  assign x392_x13_1_io_b = x391_x14_1_io_result; // @[Math.scala 152:17:@28706.4]
  assign x392_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28707.4]
  assign RetimeWrapper_60_clock = clock; // @[:@28713.4]
  assign RetimeWrapper_60_reset = reset; // @[:@28714.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28716.4]
  assign RetimeWrapper_60_io_in = x385_1_io_result; // @[package.scala 94:16:@28715.4]
  assign x393_sum_1_clock = clock; // @[:@28722.4]
  assign x393_sum_1_reset = reset; // @[:@28723.4]
  assign x393_sum_1_io_a = x392_x13_1_io_result; // @[Math.scala 151:17:@28724.4]
  assign x393_sum_1_io_b = RetimeWrapper_60_io_out; // @[Math.scala 152:17:@28725.4]
  assign x393_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28726.4]
  assign x394_1_io_b = x393_sum_1_io_result; // @[Math.scala 721:17:@28734.4]
  assign x395_mul_1_clock = clock; // @[:@28743.4]
  assign x395_mul_1_io_a = x394_1_io_result; // @[Math.scala 263:17:@28745.4]
  assign x395_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@28746.4]
  assign x395_mul_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28747.4]
  assign x396_1_io_b = x395_mul_1_io_result; // @[Math.scala 721:17:@28755.4]
  assign RetimeWrapper_61_clock = clock; // @[:@28762.4]
  assign RetimeWrapper_61_reset = reset; // @[:@28763.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28765.4]
  assign RetimeWrapper_61_io_in = x278_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@28764.4]
  assign x397_sub_1_clock = clock; // @[:@28771.4]
  assign x397_sub_1_reset = reset; // @[:@28772.4]
  assign x397_sub_1_io_a = RetimeWrapper_61_io_out; // @[Math.scala 192:17:@28773.4]
  assign x397_sub_1_io_b = x396_1_io_result; // @[Math.scala 193:17:@28774.4]
  assign x397_sub_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@28775.4]
  assign RetimeWrapper_62_clock = clock; // @[:@28784.4]
  assign RetimeWrapper_62_reset = reset; // @[:@28785.4]
  assign RetimeWrapper_62_io_flow = io_in_x242_TREADY; // @[package.scala 95:18:@28787.4]
  assign RetimeWrapper_62_io_in = 32'hf < x397_sub_number; // @[package.scala 94:16:@28786.4]
  assign x399_sub_1_clock = clock; // @[:@28793.4]
  assign x399_sub_1_reset = reset; // @[:@28794.4]
  assign x399_sub_1_io_a = x396_1_io_result; // @[Math.scala 192:17:@28795.4]
  assign x399_sub_1_io_b = RetimeWrapper_61_io_out; // @[Math.scala 193:17:@28796.4]
  assign x399_sub_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@28797.4]
  assign RetimeWrapper_63_clock = clock; // @[:@28806.4]
  assign RetimeWrapper_63_reset = reset; // @[:@28807.4]
  assign RetimeWrapper_63_io_flow = io_in_x242_TREADY; // @[package.scala 95:18:@28809.4]
  assign RetimeWrapper_63_io_in = 32'hf < x399_sub_number; // @[package.scala 94:16:@28808.4]
  assign RetimeWrapper_64_clock = clock; // @[:@28818.4]
  assign RetimeWrapper_64_reset = reset; // @[:@28819.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28821.4]
  assign RetimeWrapper_64_io_in = x397_sub_1_io_result; // @[package.scala 94:16:@28820.4]
  assign x403_1_io_b = x401 ? x571_x397_sub_D1_number : 32'h0; // @[Math.scala 721:17:@28834.4]
  assign x404_mul_1_clock = clock; // @[:@28843.4]
  assign x404_mul_1_io_a = x403_1_io_result; // @[Math.scala 263:17:@28845.4]
  assign x404_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@28846.4]
  assign x404_mul_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28847.4]
  assign x405_1_io_b = x404_mul_1_io_result; // @[Math.scala 721:17:@28855.4]
  assign RetimeWrapper_65_clock = clock; // @[:@28862.4]
  assign RetimeWrapper_65_reset = reset; // @[:@28863.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28865.4]
  assign RetimeWrapper_65_io_in = x278_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@28864.4]
  assign x406_sum_1_clock = clock; // @[:@28871.4]
  assign x406_sum_1_reset = reset; // @[:@28872.4]
  assign x406_sum_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@28873.4]
  assign x406_sum_1_io_b = x405_1_io_result; // @[Math.scala 152:17:@28874.4]
  assign x406_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28875.4]
  assign x407_1_clock = clock; // @[:@28883.4]
  assign x407_1_io_a = x278_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@28885.4]
  assign x407_1_io_b = 32'h1; // @[Math.scala 264:17:@28886.4]
  assign x407_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28887.4]
  assign x408_1_clock = clock; // @[:@28895.4]
  assign x408_1_io_a = x278_lb_0_io_rPort_9_output_0; // @[Math.scala 263:17:@28897.4]
  assign x408_1_io_b = 32'h2; // @[Math.scala 264:17:@28898.4]
  assign x408_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28899.4]
  assign x409_1_clock = clock; // @[:@28907.4]
  assign x409_1_io_a = x278_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@28909.4]
  assign x409_1_io_b = 32'h1; // @[Math.scala 264:17:@28910.4]
  assign x409_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28911.4]
  assign x410_1_clock = clock; // @[:@28919.4]
  assign x410_1_io_a = x278_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@28921.4]
  assign x410_1_io_b = 32'h2; // @[Math.scala 264:17:@28922.4]
  assign x410_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28923.4]
  assign x411_1_clock = clock; // @[:@28931.4]
  assign x411_1_io_a = x278_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@28933.4]
  assign x411_1_io_b = 32'h4; // @[Math.scala 264:17:@28934.4]
  assign x411_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28935.4]
  assign x412_1_clock = clock; // @[:@28943.4]
  assign x412_1_io_a = x278_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@28945.4]
  assign x412_1_io_b = 32'h2; // @[Math.scala 264:17:@28946.4]
  assign x412_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28947.4]
  assign x413_1_clock = clock; // @[:@28955.4]
  assign x413_1_io_a = x278_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@28957.4]
  assign x413_1_io_b = 32'h1; // @[Math.scala 264:17:@28958.4]
  assign x413_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28959.4]
  assign x414_1_clock = clock; // @[:@28967.4]
  assign x414_1_io_a = x278_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@28969.4]
  assign x414_1_io_b = 32'h2; // @[Math.scala 264:17:@28970.4]
  assign x414_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28971.4]
  assign x415_1_clock = clock; // @[:@28979.4]
  assign x415_1_io_a = x278_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@28981.4]
  assign x415_1_io_b = 32'h1; // @[Math.scala 264:17:@28982.4]
  assign x415_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@28983.4]
  assign x416_x13_1_clock = clock; // @[:@28991.4]
  assign x416_x13_1_reset = reset; // @[:@28992.4]
  assign x416_x13_1_io_a = x407_1_io_result; // @[Math.scala 151:17:@28993.4]
  assign x416_x13_1_io_b = x408_1_io_result; // @[Math.scala 152:17:@28994.4]
  assign x416_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@28995.4]
  assign x417_x14_1_clock = clock; // @[:@29001.4]
  assign x417_x14_1_reset = reset; // @[:@29002.4]
  assign x417_x14_1_io_a = x409_1_io_result; // @[Math.scala 151:17:@29003.4]
  assign x417_x14_1_io_b = x410_1_io_result; // @[Math.scala 152:17:@29004.4]
  assign x417_x14_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29005.4]
  assign x418_x13_1_clock = clock; // @[:@29011.4]
  assign x418_x13_1_reset = reset; // @[:@29012.4]
  assign x418_x13_1_io_a = x411_1_io_result; // @[Math.scala 151:17:@29013.4]
  assign x418_x13_1_io_b = x412_1_io_result; // @[Math.scala 152:17:@29014.4]
  assign x418_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29015.4]
  assign x419_x14_1_clock = clock; // @[:@29021.4]
  assign x419_x14_1_reset = reset; // @[:@29022.4]
  assign x419_x14_1_io_a = x413_1_io_result; // @[Math.scala 151:17:@29023.4]
  assign x419_x14_1_io_b = x414_1_io_result; // @[Math.scala 152:17:@29024.4]
  assign x419_x14_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29025.4]
  assign x420_x13_1_clock = clock; // @[:@29031.4]
  assign x420_x13_1_reset = reset; // @[:@29032.4]
  assign x420_x13_1_io_a = x416_x13_1_io_result; // @[Math.scala 151:17:@29033.4]
  assign x420_x13_1_io_b = x417_x14_1_io_result; // @[Math.scala 152:17:@29034.4]
  assign x420_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29035.4]
  assign x421_x14_1_clock = clock; // @[:@29041.4]
  assign x421_x14_1_reset = reset; // @[:@29042.4]
  assign x421_x14_1_io_a = x418_x13_1_io_result; // @[Math.scala 151:17:@29043.4]
  assign x421_x14_1_io_b = x419_x14_1_io_result; // @[Math.scala 152:17:@29044.4]
  assign x421_x14_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29045.4]
  assign x422_x13_1_clock = clock; // @[:@29051.4]
  assign x422_x13_1_reset = reset; // @[:@29052.4]
  assign x422_x13_1_io_a = x420_x13_1_io_result; // @[Math.scala 151:17:@29053.4]
  assign x422_x13_1_io_b = x421_x14_1_io_result; // @[Math.scala 152:17:@29054.4]
  assign x422_x13_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29055.4]
  assign RetimeWrapper_66_clock = clock; // @[:@29061.4]
  assign RetimeWrapper_66_reset = reset; // @[:@29062.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29064.4]
  assign RetimeWrapper_66_io_in = x415_1_io_result; // @[package.scala 94:16:@29063.4]
  assign x423_sum_1_clock = clock; // @[:@29070.4]
  assign x423_sum_1_reset = reset; // @[:@29071.4]
  assign x423_sum_1_io_a = x422_x13_1_io_result; // @[Math.scala 151:17:@29072.4]
  assign x423_sum_1_io_b = RetimeWrapper_66_io_out; // @[Math.scala 152:17:@29073.4]
  assign x423_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29074.4]
  assign x424_1_io_b = x423_sum_1_io_result; // @[Math.scala 721:17:@29082.4]
  assign x425_mul_1_clock = clock; // @[:@29091.4]
  assign x425_mul_1_io_a = x424_1_io_result; // @[Math.scala 263:17:@29093.4]
  assign x425_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@29094.4]
  assign x425_mul_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@29095.4]
  assign x426_1_io_b = x425_mul_1_io_result; // @[Math.scala 721:17:@29103.4]
  assign RetimeWrapper_67_clock = clock; // @[:@29110.4]
  assign RetimeWrapper_67_reset = reset; // @[:@29111.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29113.4]
  assign RetimeWrapper_67_io_in = x278_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@29112.4]
  assign x427_sub_1_clock = clock; // @[:@29119.4]
  assign x427_sub_1_reset = reset; // @[:@29120.4]
  assign x427_sub_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 192:17:@29121.4]
  assign x427_sub_1_io_b = x426_1_io_result; // @[Math.scala 193:17:@29122.4]
  assign x427_sub_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@29123.4]
  assign RetimeWrapper_68_clock = clock; // @[:@29132.4]
  assign RetimeWrapper_68_reset = reset; // @[:@29133.4]
  assign RetimeWrapper_68_io_flow = io_in_x242_TREADY; // @[package.scala 95:18:@29135.4]
  assign RetimeWrapper_68_io_in = 32'hf < x427_sub_number; // @[package.scala 94:16:@29134.4]
  assign x429_sub_1_clock = clock; // @[:@29141.4]
  assign x429_sub_1_reset = reset; // @[:@29142.4]
  assign x429_sub_1_io_a = x426_1_io_result; // @[Math.scala 192:17:@29143.4]
  assign x429_sub_1_io_b = RetimeWrapper_67_io_out; // @[Math.scala 193:17:@29144.4]
  assign x429_sub_1_io_flow = io_in_x242_TREADY; // @[Math.scala 194:20:@29145.4]
  assign RetimeWrapper_69_clock = clock; // @[:@29154.4]
  assign RetimeWrapper_69_reset = reset; // @[:@29155.4]
  assign RetimeWrapper_69_io_flow = io_in_x242_TREADY; // @[package.scala 95:18:@29157.4]
  assign RetimeWrapper_69_io_in = 32'hf < x429_sub_number; // @[package.scala 94:16:@29156.4]
  assign RetimeWrapper_70_clock = clock; // @[:@29166.4]
  assign RetimeWrapper_70_reset = reset; // @[:@29167.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29169.4]
  assign RetimeWrapper_70_io_in = x427_sub_1_io_result; // @[package.scala 94:16:@29168.4]
  assign x433_1_io_b = x431 ? x575_x427_sub_D1_number : 32'h0; // @[Math.scala 721:17:@29182.4]
  assign x434_mul_1_clock = clock; // @[:@29191.4]
  assign x434_mul_1_io_a = x433_1_io_result; // @[Math.scala 263:17:@29193.4]
  assign x434_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@29194.4]
  assign x434_mul_1_io_flow = io_in_x242_TREADY; // @[Math.scala 265:20:@29195.4]
  assign x435_1_io_b = x434_mul_1_io_result; // @[Math.scala 721:17:@29203.4]
  assign RetimeWrapper_71_clock = clock; // @[:@29210.4]
  assign RetimeWrapper_71_reset = reset; // @[:@29211.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29213.4]
  assign RetimeWrapper_71_io_in = x278_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@29212.4]
  assign x436_sum_1_clock = clock; // @[:@29219.4]
  assign x436_sum_1_reset = reset; // @[:@29220.4]
  assign x436_sum_1_io_a = RetimeWrapper_71_io_out; // @[Math.scala 151:17:@29221.4]
  assign x436_sum_1_io_b = x435_1_io_result; // @[Math.scala 152:17:@29222.4]
  assign x436_sum_1_io_flow = io_in_x242_TREADY; // @[Math.scala 153:20:@29223.4]
  assign RetimeWrapper_72_clock = clock; // @[:@29235.4]
  assign RetimeWrapper_72_reset = reset; // @[:@29236.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29238.4]
  assign RetimeWrapper_72_io_in = {x406_sum_number,x436_sum_number}; // @[package.scala 94:16:@29237.4]
  assign RetimeWrapper_73_clock = clock; // @[:@29244.4]
  assign RetimeWrapper_73_reset = reset; // @[:@29245.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29247.4]
  assign RetimeWrapper_73_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@29246.4]
  assign RetimeWrapper_74_clock = clock; // @[:@29253.4]
  assign RetimeWrapper_74_reset = reset; // @[:@29254.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29256.4]
  assign RetimeWrapper_74_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@29255.4]
  assign RetimeWrapper_75_clock = clock; // @[:@29262.4]
  assign RetimeWrapper_75_reset = reset; // @[:@29263.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29265.4]
  assign RetimeWrapper_75_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29264.4]
endmodule
module x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1( // @[:@29283.2]
  input          clock, // @[:@29284.4]
  input          reset, // @[:@29285.4]
  input          io_in_x241_TVALID, // @[:@29286.4]
  output         io_in_x241_TREADY, // @[:@29286.4]
  input  [255:0] io_in_x241_TDATA, // @[:@29286.4]
  input  [7:0]   io_in_x241_TID, // @[:@29286.4]
  input  [7:0]   io_in_x241_TDEST, // @[:@29286.4]
  output         io_in_x242_TVALID, // @[:@29286.4]
  input          io_in_x242_TREADY, // @[:@29286.4]
  output [255:0] io_in_x242_TDATA, // @[:@29286.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@29286.4]
  input          io_sigsIn_smChildAcks_0, // @[:@29286.4]
  output         io_sigsOut_smDoneIn_0, // @[:@29286.4]
  input          io_rr // @[:@29286.4]
);
  wire  x271_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire  x271_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire  x271_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire  x271_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire [12:0] x271_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire [12:0] x271_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire  x271_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire  x271_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire  x271_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@29320.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29408.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29408.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29408.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29408.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29408.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29450.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29450.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29450.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29450.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29450.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29458.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29458.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29458.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29458.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29458.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TREADY; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire [255:0] x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TDATA; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire [7:0] x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TID; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire [7:0] x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TDEST; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TVALID; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TREADY; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire [255:0] x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TDATA; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire [31:0] x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire [31:0] x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
  wire  _T_240; // @[package.scala 96:25:@29413.4 package.scala 96:25:@29414.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x442_outr_UnitPipe.scala 69:66:@29419.4]
  wire  _T_253; // @[package.scala 96:25:@29455.4 package.scala 96:25:@29456.4]
  wire  _T_259; // @[package.scala 96:25:@29463.4 package.scala 96:25:@29464.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@29466.4]
  wire  x441_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@29467.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@29475.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@29476.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@29488.4]
  x249_ctrchain x271_ctrchain ( // @[SpatialBlocks.scala 37:22:@29320.4]
    .clock(x271_ctrchain_clock),
    .reset(x271_ctrchain_reset),
    .io_input_reset(x271_ctrchain_io_input_reset),
    .io_input_enable(x271_ctrchain_io_input_enable),
    .io_output_counts_1(x271_ctrchain_io_output_counts_1),
    .io_output_counts_0(x271_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x271_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x271_ctrchain_io_output_oobs_1),
    .io_output_done(x271_ctrchain_io_output_done)
  );
  x441_inr_Foreach_SAMPLER_BOX_sm x441_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 32:18:@29380.4]
    .clock(x441_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x441_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x441_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x441_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x441_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x441_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x441_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x441_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x441_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29408.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29450.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29458.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1 x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 606:24:@29492.4]
    .clock(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x241_TREADY(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TREADY),
    .io_in_x241_TDATA(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TDATA),
    .io_in_x241_TID(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TID),
    .io_in_x241_TDEST(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TDEST),
    .io_in_x242_TVALID(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TVALID),
    .io_in_x242_TREADY(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TREADY),
    .io_in_x242_TDATA(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TDATA),
    .io_sigsIn_backpressure(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@29413.4 package.scala 96:25:@29414.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x241_TVALID | x441_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x442_outr_UnitPipe.scala 69:66:@29419.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29455.4 package.scala 96:25:@29456.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@29463.4 package.scala 96:25:@29464.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@29466.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@29467.4]
  assign _T_264 = x441_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@29475.4]
  assign _T_265 = ~ x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@29476.4]
  assign _T_272 = x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@29488.4]
  assign io_in_x241_TREADY = x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TREADY; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 48:23:@29550.4]
  assign io_in_x242_TVALID = x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TVALID; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 49:23:@29560.4]
  assign io_in_x242_TDATA = x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TDATA; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 49:23:@29558.4]
  assign io_sigsOut_smDoneIn_0 = x441_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@29473.4]
  assign x271_ctrchain_clock = clock; // @[:@29321.4]
  assign x271_ctrchain_reset = reset; // @[:@29322.4]
  assign x271_ctrchain_io_input_reset = x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@29491.4]
  assign x271_ctrchain_io_input_enable = _T_272 & x441_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@29443.4 SpatialBlocks.scala 159:42:@29490.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@29381.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@29382.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sm_io_enable = x441_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x441_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@29470.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x442_outr_UnitPipe.scala 67:50:@29416.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@29472.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x242_TREADY | x441_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@29444.4]
  assign x441_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x442_outr_UnitPipe.scala 71:48:@29422.4]
  assign RetimeWrapper_clock = clock; // @[:@29409.4]
  assign RetimeWrapper_reset = reset; // @[:@29410.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29412.4]
  assign RetimeWrapper_io_in = x271_ctrchain_io_output_done; // @[package.scala 94:16:@29411.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29451.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29452.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29454.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@29453.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29459.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29460.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29462.4]
  assign RetimeWrapper_2_io_in = x441_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@29461.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@29493.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@29494.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TDATA = io_in_x241_TDATA; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 48:23:@29549.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TID = io_in_x241_TID; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 48:23:@29545.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x241_TDEST = io_in_x241_TDEST; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 48:23:@29544.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x242_TREADY = io_in_x242_TREADY; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 49:23:@29559.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x242_TREADY | x441_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 611:22:@29577.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 611:22:@29575.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x441_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 611:22:@29573.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x271_ctrchain_io_output_counts_1[12]}},x271_ctrchain_io_output_counts_1}; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 611:22:@29568.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x271_ctrchain_io_output_counts_0[12]}},x271_ctrchain_io_output_counts_0}; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 611:22:@29567.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x271_ctrchain_io_output_oobs_0; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 611:22:@29565.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x271_ctrchain_io_output_oobs_1; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 611:22:@29566.4]
  assign x441_inr_Foreach_SAMPLER_BOX_kernelx441_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x441_inr_Foreach_SAMPLER_BOX.scala 610:18:@29561.4]
endmodule
module x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1( // @[:@29591.2]
  input          clock, // @[:@29592.4]
  input          reset, // @[:@29593.4]
  input          io_in_x241_TVALID, // @[:@29594.4]
  output         io_in_x241_TREADY, // @[:@29594.4]
  input  [255:0] io_in_x241_TDATA, // @[:@29594.4]
  input  [7:0]   io_in_x241_TID, // @[:@29594.4]
  input  [7:0]   io_in_x241_TDEST, // @[:@29594.4]
  output         io_in_x242_TVALID, // @[:@29594.4]
  input          io_in_x242_TREADY, // @[:@29594.4]
  output [255:0] io_in_x242_TDATA, // @[:@29594.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@29594.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@29594.4]
  input          io_sigsIn_smChildAcks_0, // @[:@29594.4]
  input          io_sigsIn_smChildAcks_1, // @[:@29594.4]
  output         io_sigsOut_smDoneIn_0, // @[:@29594.4]
  output         io_sigsOut_smDoneIn_1, // @[:@29594.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@29594.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@29594.4]
  input          io_rr // @[:@29594.4]
);
  wire  x244_fifoinraw_0_clock; // @[m_x244_fifoinraw_0.scala 27:17:@29608.4]
  wire  x244_fifoinraw_0_reset; // @[m_x244_fifoinraw_0.scala 27:17:@29608.4]
  wire  x245_fifoinpacked_0_clock; // @[m_x245_fifoinpacked_0.scala 27:17:@29632.4]
  wire  x245_fifoinpacked_0_reset; // @[m_x245_fifoinpacked_0.scala 27:17:@29632.4]
  wire  x245_fifoinpacked_0_io_wPort_0_en_0; // @[m_x245_fifoinpacked_0.scala 27:17:@29632.4]
  wire  x245_fifoinpacked_0_io_full; // @[m_x245_fifoinpacked_0.scala 27:17:@29632.4]
  wire  x245_fifoinpacked_0_io_active_0_in; // @[m_x245_fifoinpacked_0.scala 27:17:@29632.4]
  wire  x245_fifoinpacked_0_io_active_0_out; // @[m_x245_fifoinpacked_0.scala 27:17:@29632.4]
  wire  x246_fifooutraw_0_clock; // @[m_x246_fifooutraw_0.scala 27:17:@29656.4]
  wire  x246_fifooutraw_0_reset; // @[m_x246_fifooutraw_0.scala 27:17:@29656.4]
  wire  x249_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire  x249_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire  x249_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire  x249_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire [12:0] x249_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire [12:0] x249_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire  x249_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire  x249_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire  x249_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@29680.4]
  wire  x267_inr_Foreach_sm_clock; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_reset; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_enable; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_done; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_doneLatch; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_ctrDone; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_datapathEn; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_ctrInc; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_ctrRst; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_parentAck; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_backpressure; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  x267_inr_Foreach_sm_io_break; // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29768.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29768.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29768.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29768.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29768.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29814.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29814.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29814.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29814.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29814.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29822.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29822.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29822.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29822.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29822.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_clock; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_reset; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_wPort_0_en_0; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_full; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_active_0_in; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_active_0_out; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire [31:0] x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire [31:0] x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_rr; // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
  wire  x442_outr_UnitPipe_sm_clock; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_reset; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_enable; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_done; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_rst; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_ctrDone; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_ctrInc; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_parentAck; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  x442_outr_UnitPipe_sm_io_childAck_0; // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30046.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30046.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30046.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30046.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30046.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30054.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30054.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30054.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30054.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30054.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_clock; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_reset; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TVALID; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TREADY; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire [255:0] x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TDATA; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire [7:0] x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TID; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire [7:0] x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TDEST; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TVALID; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TREADY; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire [255:0] x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TDATA; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_rr; // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
  wire  _T_254; // @[package.scala 96:25:@29773.4 package.scala 96:25:@29774.4]
  wire  _T_260; // @[implicits.scala 47:10:@29777.4]
  wire  _T_261; // @[sm_x443_outr_UnitPipe.scala 70:41:@29778.4]
  wire  _T_262; // @[sm_x443_outr_UnitPipe.scala 70:78:@29779.4]
  wire  _T_263; // @[sm_x443_outr_UnitPipe.scala 70:76:@29780.4]
  wire  _T_275; // @[package.scala 96:25:@29819.4 package.scala 96:25:@29820.4]
  wire  _T_281; // @[package.scala 96:25:@29827.4 package.scala 96:25:@29828.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@29830.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@29839.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@29840.4]
  wire  _T_354; // @[package.scala 100:49:@30017.4]
  reg  _T_357; // @[package.scala 48:56:@30018.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@30051.4 package.scala 96:25:@30052.4]
  wire  _T_377; // @[package.scala 96:25:@30059.4 package.scala 96:25:@30060.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@30062.4]
  x244_fifoinraw_0 x244_fifoinraw_0 ( // @[m_x244_fifoinraw_0.scala 27:17:@29608.4]
    .clock(x244_fifoinraw_0_clock),
    .reset(x244_fifoinraw_0_reset)
  );
  x245_fifoinpacked_0 x245_fifoinpacked_0 ( // @[m_x245_fifoinpacked_0.scala 27:17:@29632.4]
    .clock(x245_fifoinpacked_0_clock),
    .reset(x245_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x245_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x245_fifoinpacked_0_io_full),
    .io_active_0_in(x245_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x245_fifoinpacked_0_io_active_0_out)
  );
  x244_fifoinraw_0 x246_fifooutraw_0 ( // @[m_x246_fifooutraw_0.scala 27:17:@29656.4]
    .clock(x246_fifooutraw_0_clock),
    .reset(x246_fifooutraw_0_reset)
  );
  x249_ctrchain x249_ctrchain ( // @[SpatialBlocks.scala 37:22:@29680.4]
    .clock(x249_ctrchain_clock),
    .reset(x249_ctrchain_reset),
    .io_input_reset(x249_ctrchain_io_input_reset),
    .io_input_enable(x249_ctrchain_io_input_enable),
    .io_output_counts_1(x249_ctrchain_io_output_counts_1),
    .io_output_counts_0(x249_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x249_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x249_ctrchain_io_output_oobs_1),
    .io_output_done(x249_ctrchain_io_output_done)
  );
  x267_inr_Foreach_sm x267_inr_Foreach_sm ( // @[sm_x267_inr_Foreach.scala 32:18:@29740.4]
    .clock(x267_inr_Foreach_sm_clock),
    .reset(x267_inr_Foreach_sm_reset),
    .io_enable(x267_inr_Foreach_sm_io_enable),
    .io_done(x267_inr_Foreach_sm_io_done),
    .io_doneLatch(x267_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x267_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x267_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x267_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x267_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x267_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x267_inr_Foreach_sm_io_backpressure),
    .io_break(x267_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29768.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29814.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29822.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x267_inr_Foreach_kernelx267_inr_Foreach_concrete1 x267_inr_Foreach_kernelx267_inr_Foreach_concrete1 ( // @[sm_x267_inr_Foreach.scala 106:24:@29857.4]
    .clock(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_clock),
    .reset(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_reset),
    .io_in_x245_fifoinpacked_0_wPort_0_en_0(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_wPort_0_en_0),
    .io_in_x245_fifoinpacked_0_full(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_full),
    .io_in_x245_fifoinpacked_0_active_0_in(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_active_0_in),
    .io_in_x245_fifoinpacked_0_active_0_out(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x442_outr_UnitPipe_sm ( // @[sm_x442_outr_UnitPipe.scala 32:18:@29989.4]
    .clock(x442_outr_UnitPipe_sm_clock),
    .reset(x442_outr_UnitPipe_sm_reset),
    .io_enable(x442_outr_UnitPipe_sm_io_enable),
    .io_done(x442_outr_UnitPipe_sm_io_done),
    .io_rst(x442_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x442_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x442_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x442_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x442_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x442_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x442_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30046.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30054.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1 x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1 ( // @[sm_x442_outr_UnitPipe.scala 76:24:@30084.4]
    .clock(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_clock),
    .reset(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_reset),
    .io_in_x241_TVALID(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TVALID),
    .io_in_x241_TREADY(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TREADY),
    .io_in_x241_TDATA(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TDATA),
    .io_in_x241_TID(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TID),
    .io_in_x241_TDEST(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TDEST),
    .io_in_x242_TVALID(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TVALID),
    .io_in_x242_TREADY(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TREADY),
    .io_in_x242_TDATA(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TDATA),
    .io_sigsIn_smEnableOuts_0(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@29773.4 package.scala 96:25:@29774.4]
  assign _T_260 = x245_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@29777.4]
  assign _T_261 = ~ _T_260; // @[sm_x443_outr_UnitPipe.scala 70:41:@29778.4]
  assign _T_262 = ~ x245_fifoinpacked_0_io_active_0_out; // @[sm_x443_outr_UnitPipe.scala 70:78:@29779.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x443_outr_UnitPipe.scala 70:76:@29780.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29819.4 package.scala 96:25:@29820.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@29827.4 package.scala 96:25:@29828.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@29830.4]
  assign _T_286 = x267_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@29839.4]
  assign _T_287 = ~ x267_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@29840.4]
  assign _T_354 = x442_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@30017.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30051.4 package.scala 96:25:@30052.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30059.4 package.scala 96:25:@30060.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@30062.4]
  assign io_in_x241_TREADY = x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TREADY; // @[sm_x442_outr_UnitPipe.scala 48:23:@30140.4]
  assign io_in_x242_TVALID = x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TVALID; // @[sm_x442_outr_UnitPipe.scala 49:23:@30150.4]
  assign io_in_x242_TDATA = x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TDATA; // @[sm_x442_outr_UnitPipe.scala 49:23:@30148.4]
  assign io_sigsOut_smDoneIn_0 = x267_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@29837.4]
  assign io_sigsOut_smDoneIn_1 = x442_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@30069.4]
  assign io_sigsOut_smCtrCopyDone_0 = x267_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@29856.4]
  assign io_sigsOut_smCtrCopyDone_1 = x442_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@30083.4]
  assign x244_fifoinraw_0_clock = clock; // @[:@29609.4]
  assign x244_fifoinraw_0_reset = reset; // @[:@29610.4]
  assign x245_fifoinpacked_0_clock = clock; // @[:@29633.4]
  assign x245_fifoinpacked_0_reset = reset; // @[:@29634.4]
  assign x245_fifoinpacked_0_io_wPort_0_en_0 = x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@29917.4]
  assign x245_fifoinpacked_0_io_active_0_in = x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@29916.4]
  assign x246_fifooutraw_0_clock = clock; // @[:@29657.4]
  assign x246_fifooutraw_0_reset = reset; // @[:@29658.4]
  assign x249_ctrchain_clock = clock; // @[:@29681.4]
  assign x249_ctrchain_reset = reset; // @[:@29682.4]
  assign x249_ctrchain_io_input_reset = x267_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@29855.4]
  assign x249_ctrchain_io_input_enable = x267_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@29807.4 SpatialBlocks.scala 159:42:@29854.4]
  assign x267_inr_Foreach_sm_clock = clock; // @[:@29741.4]
  assign x267_inr_Foreach_sm_reset = reset; // @[:@29742.4]
  assign x267_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@29834.4]
  assign x267_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x443_outr_UnitPipe.scala 69:38:@29776.4]
  assign x267_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@29836.4]
  assign x267_inr_Foreach_sm_io_backpressure = _T_263 | x267_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@29808.4]
  assign x267_inr_Foreach_sm_io_break = 1'h0; // @[sm_x443_outr_UnitPipe.scala 73:36:@29786.4]
  assign RetimeWrapper_clock = clock; // @[:@29769.4]
  assign RetimeWrapper_reset = reset; // @[:@29770.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29772.4]
  assign RetimeWrapper_io_in = x249_ctrchain_io_output_done; // @[package.scala 94:16:@29771.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29815.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29816.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29818.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@29817.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29823.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29824.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29826.4]
  assign RetimeWrapper_2_io_in = x267_inr_Foreach_sm_io_done; // @[package.scala 94:16:@29825.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_clock = clock; // @[:@29858.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_reset = reset; // @[:@29859.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_full = x245_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@29911.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_in_x245_fifoinpacked_0_active_0_out = x245_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@29910.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x267_inr_Foreach_sm_io_doneLatch; // @[sm_x267_inr_Foreach.scala 111:22:@29940.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x267_inr_Foreach.scala 111:22:@29938.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_break = x267_inr_Foreach_sm_io_break; // @[sm_x267_inr_Foreach.scala 111:22:@29936.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x249_ctrchain_io_output_counts_1[12]}},x249_ctrchain_io_output_counts_1}; // @[sm_x267_inr_Foreach.scala 111:22:@29931.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x249_ctrchain_io_output_counts_0[12]}},x249_ctrchain_io_output_counts_0}; // @[sm_x267_inr_Foreach.scala 111:22:@29930.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x249_ctrchain_io_output_oobs_0; // @[sm_x267_inr_Foreach.scala 111:22:@29928.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x249_ctrchain_io_output_oobs_1; // @[sm_x267_inr_Foreach.scala 111:22:@29929.4]
  assign x267_inr_Foreach_kernelx267_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x267_inr_Foreach.scala 110:18:@29924.4]
  assign x442_outr_UnitPipe_sm_clock = clock; // @[:@29990.4]
  assign x442_outr_UnitPipe_sm_reset = reset; // @[:@29991.4]
  assign x442_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@30066.4]
  assign x442_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@30041.4]
  assign x442_outr_UnitPipe_sm_io_ctrDone = x442_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x443_outr_UnitPipe.scala 78:40:@30021.4]
  assign x442_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@30068.4]
  assign x442_outr_UnitPipe_sm_io_doneIn_0 = x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@30038.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30047.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30048.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30050.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@30049.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30055.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30056.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30058.4]
  assign RetimeWrapper_4_io_in = x442_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@30057.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_clock = clock; // @[:@30085.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_reset = reset; // @[:@30086.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TVALID = io_in_x241_TVALID; // @[sm_x442_outr_UnitPipe.scala 48:23:@30141.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TDATA = io_in_x241_TDATA; // @[sm_x442_outr_UnitPipe.scala 48:23:@30139.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TID = io_in_x241_TID; // @[sm_x442_outr_UnitPipe.scala 48:23:@30135.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x241_TDEST = io_in_x241_TDEST; // @[sm_x442_outr_UnitPipe.scala 48:23:@30134.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_in_x242_TREADY = io_in_x242_TREADY; // @[sm_x442_outr_UnitPipe.scala 49:23:@30149.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x442_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x442_outr_UnitPipe.scala 81:22:@30159.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x442_outr_UnitPipe_sm_io_childAck_0; // @[sm_x442_outr_UnitPipe.scala 81:22:@30157.4]
  assign x442_outr_UnitPipe_kernelx442_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x442_outr_UnitPipe.scala 80:18:@30151.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x465_outr_UnitPipe_sm( // @[:@30648.2]
  input   clock, // @[:@30649.4]
  input   reset, // @[:@30650.4]
  input   io_enable, // @[:@30651.4]
  output  io_done, // @[:@30651.4]
  input   io_parentAck, // @[:@30651.4]
  input   io_doneIn_0, // @[:@30651.4]
  input   io_doneIn_1, // @[:@30651.4]
  input   io_doneIn_2, // @[:@30651.4]
  output  io_enableOut_0, // @[:@30651.4]
  output  io_enableOut_1, // @[:@30651.4]
  output  io_enableOut_2, // @[:@30651.4]
  output  io_childAck_0, // @[:@30651.4]
  output  io_childAck_1, // @[:@30651.4]
  output  io_childAck_2, // @[:@30651.4]
  input   io_ctrCopyDone_0, // @[:@30651.4]
  input   io_ctrCopyDone_1, // @[:@30651.4]
  input   io_ctrCopyDone_2 // @[:@30651.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@30654.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@30654.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@30654.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@30654.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@30654.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@30654.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@30657.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@30657.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@30657.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@30657.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@30657.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@30657.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@30660.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@30660.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@30660.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@30660.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@30660.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@30660.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@30663.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@30663.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@30663.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@30663.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@30663.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@30663.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@30666.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@30666.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@30666.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@30666.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@30666.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@30666.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@30669.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@30669.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@30669.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@30669.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@30669.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@30669.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@30710.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@30710.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@30710.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@30710.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@30710.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@30710.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@30713.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@30713.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@30713.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@30713.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@30713.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@30713.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@30716.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@30716.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@30716.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@30716.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@30716.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@30716.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30767.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30767.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30767.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30767.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30767.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30781.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30781.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30781.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30781.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30781.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30836.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30836.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30836.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30836.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30836.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30850.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30850.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30850.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30850.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30850.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@30868.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@30868.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@30868.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@30868.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@30868.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@30905.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@30905.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@30905.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@30905.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@30905.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@30919.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@30919.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@30919.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@30919.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@30919.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@30937.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@30937.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@30937.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@30937.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@30937.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@30994.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@30994.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@30994.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@30994.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@30994.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@31011.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@31011.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@31011.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@31011.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@31011.4]
  wire  _T_77; // @[Controllers.scala 80:47:@30672.4]
  wire  allDone; // @[Controllers.scala 80:47:@30673.4]
  wire  _T_151; // @[Controllers.scala 165:35:@30751.4]
  wire  _T_153; // @[Controllers.scala 165:60:@30752.4]
  wire  _T_154; // @[Controllers.scala 165:58:@30753.4]
  wire  _T_156; // @[Controllers.scala 165:76:@30754.4]
  wire  _T_157; // @[Controllers.scala 165:74:@30755.4]
  wire  _T_161; // @[Controllers.scala 165:109:@30758.4]
  wire  _T_164; // @[Controllers.scala 165:141:@30760.4]
  wire  _T_172; // @[package.scala 96:25:@30772.4 package.scala 96:25:@30773.4]
  wire  _T_176; // @[Controllers.scala 167:54:@30775.4]
  wire  _T_177; // @[Controllers.scala 167:52:@30776.4]
  wire  _T_184; // @[package.scala 96:25:@30786.4 package.scala 96:25:@30787.4]
  wire  _T_202; // @[package.scala 96:25:@30804.4 package.scala 96:25:@30805.4]
  wire  _T_206; // @[Controllers.scala 169:67:@30807.4]
  wire  _T_207; // @[Controllers.scala 169:86:@30808.4]
  wire  _T_219; // @[Controllers.scala 165:35:@30820.4]
  wire  _T_221; // @[Controllers.scala 165:60:@30821.4]
  wire  _T_222; // @[Controllers.scala 165:58:@30822.4]
  wire  _T_224; // @[Controllers.scala 165:76:@30823.4]
  wire  _T_225; // @[Controllers.scala 165:74:@30824.4]
  wire  _T_229; // @[Controllers.scala 165:109:@30827.4]
  wire  _T_232; // @[Controllers.scala 165:141:@30829.4]
  wire  _T_240; // @[package.scala 96:25:@30841.4 package.scala 96:25:@30842.4]
  wire  _T_244; // @[Controllers.scala 167:54:@30844.4]
  wire  _T_245; // @[Controllers.scala 167:52:@30845.4]
  wire  _T_252; // @[package.scala 96:25:@30855.4 package.scala 96:25:@30856.4]
  wire  _T_270; // @[package.scala 96:25:@30873.4 package.scala 96:25:@30874.4]
  wire  _T_274; // @[Controllers.scala 169:67:@30876.4]
  wire  _T_275; // @[Controllers.scala 169:86:@30877.4]
  wire  _T_287; // @[Controllers.scala 165:35:@30889.4]
  wire  _T_289; // @[Controllers.scala 165:60:@30890.4]
  wire  _T_290; // @[Controllers.scala 165:58:@30891.4]
  wire  _T_292; // @[Controllers.scala 165:76:@30892.4]
  wire  _T_293; // @[Controllers.scala 165:74:@30893.4]
  wire  _T_297; // @[Controllers.scala 165:109:@30896.4]
  wire  _T_300; // @[Controllers.scala 165:141:@30898.4]
  wire  _T_308; // @[package.scala 96:25:@30910.4 package.scala 96:25:@30911.4]
  wire  _T_312; // @[Controllers.scala 167:54:@30913.4]
  wire  _T_313; // @[Controllers.scala 167:52:@30914.4]
  wire  _T_320; // @[package.scala 96:25:@30924.4 package.scala 96:25:@30925.4]
  wire  _T_338; // @[package.scala 96:25:@30942.4 package.scala 96:25:@30943.4]
  wire  _T_342; // @[Controllers.scala 169:67:@30945.4]
  wire  _T_343; // @[Controllers.scala 169:86:@30946.4]
  wire  _T_358; // @[Controllers.scala 213:68:@30964.4]
  wire  _T_360; // @[Controllers.scala 213:90:@30966.4]
  wire  _T_362; // @[Controllers.scala 213:132:@30968.4]
  wire  _T_366; // @[Controllers.scala 213:68:@30973.4]
  wire  _T_368; // @[Controllers.scala 213:90:@30975.4]
  wire  _T_374; // @[Controllers.scala 213:68:@30981.4]
  wire  _T_376; // @[Controllers.scala 213:90:@30983.4]
  wire  _T_383; // @[package.scala 100:49:@30989.4]
  reg  _T_386; // @[package.scala 48:56:@30990.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@30992.4]
  reg  _T_400; // @[package.scala 48:56:@31008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@30654.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@30657.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@30660.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@30663.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@30666.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@30669.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@30710.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@30713.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@30716.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30767.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30781.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30799.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30836.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30850.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@30868.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@30905.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@30919.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@30937.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@30994.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@31011.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@30672.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@30673.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@30751.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@30752.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@30753.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@30754.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@30755.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@30758.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@30760.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@30772.4 package.scala 96:25:@30773.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@30775.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@30776.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30786.4 package.scala 96:25:@30787.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@30804.4 package.scala 96:25:@30805.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@30807.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@30808.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@30820.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@30821.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@30822.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@30823.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@30824.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@30827.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@30829.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30841.4 package.scala 96:25:@30842.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@30844.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@30845.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30855.4 package.scala 96:25:@30856.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@30873.4 package.scala 96:25:@30874.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@30876.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@30877.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@30889.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@30890.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@30891.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@30892.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@30893.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@30896.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@30898.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@30910.4 package.scala 96:25:@30911.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@30913.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@30914.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@30924.4 package.scala 96:25:@30925.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@30942.4 package.scala 96:25:@30943.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@30945.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@30946.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@30964.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@30966.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@30968.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@30973.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@30975.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@30981.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@30983.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@30989.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@30992.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@31018.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@30972.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@30980.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@30988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@30959.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@30961.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@30963.4]
  assign active_0_clock = clock; // @[:@30655.4]
  assign active_0_reset = reset; // @[:@30656.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@30762.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@30766.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30676.4]
  assign active_1_clock = clock; // @[:@30658.4]
  assign active_1_reset = reset; // @[:@30659.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@30831.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@30835.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30677.4]
  assign active_2_clock = clock; // @[:@30661.4]
  assign active_2_reset = reset; // @[:@30662.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@30900.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@30904.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30678.4]
  assign done_0_clock = clock; // @[:@30664.4]
  assign done_0_reset = reset; // @[:@30665.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@30812.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30690.4 Controllers.scala 170:32:@30819.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30679.4]
  assign done_1_clock = clock; // @[:@30667.4]
  assign done_1_reset = reset; // @[:@30668.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@30881.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30699.4 Controllers.scala 170:32:@30888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30680.4]
  assign done_2_clock = clock; // @[:@30670.4]
  assign done_2_reset = reset; // @[:@30671.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@30950.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30708.4 Controllers.scala 170:32:@30957.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30681.4]
  assign iterDone_0_clock = clock; // @[:@30711.4]
  assign iterDone_0_reset = reset; // @[:@30712.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@30780.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@30730.4 Controllers.scala 168:36:@30796.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30719.4]
  assign iterDone_1_clock = clock; // @[:@30714.4]
  assign iterDone_1_reset = reset; // @[:@30715.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@30849.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@30739.4 Controllers.scala 168:36:@30865.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30720.4]
  assign iterDone_2_clock = clock; // @[:@30717.4]
  assign iterDone_2_reset = reset; // @[:@30718.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@30918.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@30748.4 Controllers.scala 168:36:@30934.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30721.4]
  assign RetimeWrapper_clock = clock; // @[:@30768.4]
  assign RetimeWrapper_reset = reset; // @[:@30769.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30771.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@30770.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30782.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30783.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30785.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@30784.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30800.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30801.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30803.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@30802.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30837.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30838.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30840.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@30839.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30851.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30852.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30854.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@30853.4]
  assign RetimeWrapper_5_clock = clock; // @[:@30869.4]
  assign RetimeWrapper_5_reset = reset; // @[:@30870.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@30872.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@30871.4]
  assign RetimeWrapper_6_clock = clock; // @[:@30906.4]
  assign RetimeWrapper_6_reset = reset; // @[:@30907.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@30909.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@30908.4]
  assign RetimeWrapper_7_clock = clock; // @[:@30920.4]
  assign RetimeWrapper_7_reset = reset; // @[:@30921.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@30923.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@30922.4]
  assign RetimeWrapper_8_clock = clock; // @[:@30938.4]
  assign RetimeWrapper_8_reset = reset; // @[:@30939.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@30941.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@30940.4]
  assign RetimeWrapper_9_clock = clock; // @[:@30995.4]
  assign RetimeWrapper_9_reset = reset; // @[:@30996.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@30998.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@30997.4]
  assign RetimeWrapper_10_clock = clock; // @[:@31012.4]
  assign RetimeWrapper_10_reset = reset; // @[:@31013.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@31015.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@31014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x451_inr_UnitPipe_sm( // @[:@31191.2]
  input   clock, // @[:@31192.4]
  input   reset, // @[:@31193.4]
  input   io_enable, // @[:@31194.4]
  output  io_done, // @[:@31194.4]
  output  io_doneLatch, // @[:@31194.4]
  input   io_ctrDone, // @[:@31194.4]
  output  io_datapathEn, // @[:@31194.4]
  output  io_ctrInc, // @[:@31194.4]
  input   io_parentAck, // @[:@31194.4]
  input   io_backpressure // @[:@31194.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@31196.4]
  wire  active_reset; // @[Controllers.scala 261:22:@31196.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@31196.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@31196.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@31196.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@31196.4]
  wire  done_clock; // @[Controllers.scala 262:20:@31199.4]
  wire  done_reset; // @[Controllers.scala 262:20:@31199.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@31199.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@31199.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@31199.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@31199.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31253.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31253.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31253.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31253.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31253.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31261.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31261.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31261.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31261.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31261.4]
  wire  _T_80; // @[Controllers.scala 264:48:@31204.4]
  wire  _T_81; // @[Controllers.scala 264:46:@31205.4]
  wire  _T_82; // @[Controllers.scala 264:62:@31206.4]
  wire  _T_83; // @[Controllers.scala 264:60:@31207.4]
  wire  _T_100; // @[package.scala 100:49:@31224.4]
  reg  _T_103; // @[package.scala 48:56:@31225.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@31233.4]
  wire  _T_116; // @[Controllers.scala 283:41:@31241.4]
  wire  _T_117; // @[Controllers.scala 283:59:@31242.4]
  wire  _T_119; // @[Controllers.scala 284:37:@31245.4]
  reg  _T_125; // @[package.scala 48:56:@31249.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@31271.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@31274.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@31276.4]
  wire  _T_152; // @[Controllers.scala 292:61:@31277.4]
  wire  _T_153; // @[Controllers.scala 292:24:@31278.4]
  SRFF active ( // @[Controllers.scala 261:22:@31196.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@31199.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31253.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31261.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@31204.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@31205.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@31206.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@31207.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@31224.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@31233.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@31241.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@31242.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@31245.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@31276.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@31277.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@31278.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@31252.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@31280.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@31244.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@31247.4]
  assign active_clock = clock; // @[:@31197.4]
  assign active_reset = reset; // @[:@31198.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@31209.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@31213.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@31214.4]
  assign done_clock = clock; // @[:@31200.4]
  assign done_reset = reset; // @[:@31201.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@31229.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@31222.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@31223.4]
  assign RetimeWrapper_clock = clock; // @[:@31254.4]
  assign RetimeWrapper_reset = reset; // @[:@31255.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31257.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@31256.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31262.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31263.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31265.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@31264.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1( // @[:@31355.2]
  output        io_in_x444_valid, // @[:@31358.4]
  output [63:0] io_in_x444_bits_addr, // @[:@31358.4]
  output [31:0] io_in_x444_bits_size, // @[:@31358.4]
  input  [63:0] io_in_x239_outdram_number, // @[:@31358.4]
  input         io_sigsIn_backpressure, // @[:@31358.4]
  input         io_sigsIn_datapathEn, // @[:@31358.4]
  input         io_rr // @[:@31358.4]
);
  wire [96:0] x448_tuple; // @[Cat.scala 30:58:@31372.4]
  wire  _T_135; // @[implicits.scala 55:10:@31375.4]
  assign x448_tuple = {33'h7e9000,io_in_x239_outdram_number}; // @[Cat.scala 30:58:@31372.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@31375.4]
  assign io_in_x444_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x451_inr_UnitPipe.scala 65:18:@31378.4]
  assign io_in_x444_bits_addr = x448_tuple[63:0]; // @[sm_x451_inr_UnitPipe.scala 66:22:@31380.4]
  assign io_in_x444_bits_size = x448_tuple[95:64]; // @[sm_x451_inr_UnitPipe.scala 67:22:@31382.4]
endmodule
module FF_13( // @[:@31384.2]
  input         clock, // @[:@31385.4]
  input         reset, // @[:@31386.4]
  output [22:0] io_rPort_0_output_0, // @[:@31387.4]
  input  [22:0] io_wPort_0_data_0, // @[:@31387.4]
  input         io_wPort_0_reset, // @[:@31387.4]
  input         io_wPort_0_en_0 // @[:@31387.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@31402.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@31404.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@31405.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@31404.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@31405.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@31407.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@31422.2]
  input         clock, // @[:@31423.4]
  input         reset, // @[:@31424.4]
  input         io_input_reset, // @[:@31425.4]
  input         io_input_enable, // @[:@31425.4]
  output [22:0] io_output_count_0, // @[:@31425.4]
  output        io_output_oobs_0, // @[:@31425.4]
  output        io_output_done // @[:@31425.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@31438.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@31438.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@31438.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@31438.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@31438.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@31438.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@31454.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@31454.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@31454.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@31454.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@31454.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@31454.4]
  wire  _T_36; // @[Counter.scala 264:45:@31457.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@31482.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@31483.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@31484.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@31485.4]
  wire  _T_57; // @[Counter.scala 293:18:@31487.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@31495.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@31498.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@31499.4]
  wire  _T_75; // @[Counter.scala 322:102:@31503.4]
  wire  _T_77; // @[Counter.scala 322:130:@31504.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@31438.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@31454.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@31457.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@31482.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@31483.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@31484.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@31485.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@31487.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@31495.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@31498.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@31499.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@31503.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@31504.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@31502.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@31506.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@31508.4]
  assign bases_0_clock = clock; // @[:@31439.4]
  assign bases_0_reset = reset; // @[:@31440.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@31501.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@31480.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@31481.4]
  assign SRFF_clock = clock; // @[:@31455.4]
  assign SRFF_reset = reset; // @[:@31456.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@31459.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@31461.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@31462.4]
endmodule
module x453_ctrchain( // @[:@31513.2]
  input         clock, // @[:@31514.4]
  input         reset, // @[:@31515.4]
  input         io_input_reset, // @[:@31516.4]
  input         io_input_enable, // @[:@31516.4]
  output [22:0] io_output_counts_0, // @[:@31516.4]
  output        io_output_oobs_0, // @[:@31516.4]
  output        io_output_done // @[:@31516.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@31518.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@31518.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@31518.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@31518.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@31518.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@31518.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@31518.4]
  reg  wasDone; // @[Counter.scala 542:24:@31527.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@31533.4]
  wire  _T_47; // @[Counter.scala 546:80:@31534.4]
  reg  doneLatch; // @[Counter.scala 550:26:@31539.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@31540.4]
  wire  _T_55; // @[Counter.scala 551:19:@31541.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@31518.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@31533.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@31534.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@31540.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@31541.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@31543.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@31545.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@31536.4]
  assign ctrs_0_clock = clock; // @[:@31519.4]
  assign ctrs_0_reset = reset; // @[:@31520.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@31524.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@31525.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x460_inr_Foreach_sm( // @[:@31733.2]
  input   clock, // @[:@31734.4]
  input   reset, // @[:@31735.4]
  input   io_enable, // @[:@31736.4]
  output  io_done, // @[:@31736.4]
  output  io_doneLatch, // @[:@31736.4]
  input   io_ctrDone, // @[:@31736.4]
  output  io_datapathEn, // @[:@31736.4]
  output  io_ctrInc, // @[:@31736.4]
  output  io_ctrRst, // @[:@31736.4]
  input   io_parentAck, // @[:@31736.4]
  input   io_backpressure, // @[:@31736.4]
  input   io_break // @[:@31736.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@31738.4]
  wire  active_reset; // @[Controllers.scala 261:22:@31738.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@31738.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@31738.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@31738.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@31738.4]
  wire  done_clock; // @[Controllers.scala 262:20:@31741.4]
  wire  done_reset; // @[Controllers.scala 262:20:@31741.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@31741.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@31741.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@31741.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@31741.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31775.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31775.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31775.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31775.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31775.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31797.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31797.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31797.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31797.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31797.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31817.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31817.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31817.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31817.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31817.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@31833.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@31833.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@31833.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@31833.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@31833.4]
  wire  _T_80; // @[Controllers.scala 264:48:@31746.4]
  wire  _T_81; // @[Controllers.scala 264:46:@31747.4]
  wire  _T_82; // @[Controllers.scala 264:62:@31748.4]
  wire  _T_83; // @[Controllers.scala 264:60:@31749.4]
  wire  _T_100; // @[package.scala 100:49:@31766.4]
  reg  _T_103; // @[package.scala 48:56:@31767.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@31780.4 package.scala 96:25:@31781.4]
  wire  _T_110; // @[package.scala 100:49:@31782.4]
  reg  _T_113; // @[package.scala 48:56:@31783.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@31785.4]
  wire  _T_118; // @[Controllers.scala 283:41:@31790.4]
  wire  _T_119; // @[Controllers.scala 283:59:@31791.4]
  wire  _T_121; // @[Controllers.scala 284:37:@31794.4]
  wire  _T_124; // @[package.scala 96:25:@31802.4 package.scala 96:25:@31803.4]
  wire  _T_126; // @[package.scala 100:49:@31804.4]
  reg  _T_129; // @[package.scala 48:56:@31805.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@31827.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@31829.4]
  reg  _T_153; // @[package.scala 48:56:@31830.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@31838.4 package.scala 96:25:@31839.4]
  wire  _T_158; // @[Controllers.scala 292:61:@31840.4]
  wire  _T_159; // @[Controllers.scala 292:24:@31841.4]
  SRFF active ( // @[Controllers.scala 261:22:@31738.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@31741.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@31775.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@31797.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31809.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31817.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@31833.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@31746.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@31747.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@31748.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@31749.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@31766.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@31780.4 package.scala 96:25:@31781.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@31782.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@31785.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@31790.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@31791.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@31794.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31802.4 package.scala 96:25:@31803.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@31804.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@31829.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@31838.4 package.scala 96:25:@31839.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@31840.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@31841.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@31808.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@31843.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@31793.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@31796.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@31788.4]
  assign active_clock = clock; // @[:@31739.4]
  assign active_reset = reset; // @[:@31740.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@31751.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@31755.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@31756.4]
  assign done_clock = clock; // @[:@31742.4]
  assign done_reset = reset; // @[:@31743.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@31771.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@31764.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@31765.4]
  assign RetimeWrapper_clock = clock; // @[:@31776.4]
  assign RetimeWrapper_reset = reset; // @[:@31777.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@31779.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@31778.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31798.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31799.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@31801.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@31800.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31810.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31811.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31813.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@31812.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31818.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31819.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31821.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@31820.4]
  assign RetimeWrapper_4_clock = clock; // @[:@31834.4]
  assign RetimeWrapper_4_reset = reset; // @[:@31835.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@31837.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@31836.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x460_inr_Foreach_kernelx460_inr_Foreach_concrete1( // @[:@32050.2]
  input         clock, // @[:@32051.4]
  input         reset, // @[:@32052.4]
  output [20:0] io_in_x243_outbuf_0_rPort_0_ofs_0, // @[:@32053.4]
  output        io_in_x243_outbuf_0_rPort_0_en_0, // @[:@32053.4]
  output        io_in_x243_outbuf_0_rPort_0_backpressure, // @[:@32053.4]
  input  [31:0] io_in_x243_outbuf_0_rPort_0_output_0, // @[:@32053.4]
  output        io_in_x445_valid, // @[:@32053.4]
  output [31:0] io_in_x445_bits_wdata_0, // @[:@32053.4]
  output        io_in_x445_bits_wstrb, // @[:@32053.4]
  input         io_sigsIn_backpressure, // @[:@32053.4]
  input         io_sigsIn_datapathEn, // @[:@32053.4]
  input         io_sigsIn_break, // @[:@32053.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@32053.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@32053.4]
  input         io_rr // @[:@32053.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@32080.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@32080.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32109.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32109.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32109.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32109.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32109.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32118.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32118.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32118.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32118.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32118.4]
  wire  b455; // @[sm_x460_inr_Foreach.scala 62:18:@32088.4]
  wire  _T_274; // @[sm_x460_inr_Foreach.scala 67:129:@32092.4]
  wire  _T_278; // @[implicits.scala 55:10:@32095.4]
  wire  _T_279; // @[sm_x460_inr_Foreach.scala 67:146:@32096.4]
  wire [32:0] x458_tuple; // @[Cat.scala 30:58:@32106.4]
  wire  _T_290; // @[package.scala 96:25:@32123.4 package.scala 96:25:@32124.4]
  wire  _T_292; // @[implicits.scala 55:10:@32125.4]
  wire  x579_b455_D2; // @[package.scala 96:25:@32114.4 package.scala 96:25:@32115.4]
  wire  _T_293; // @[sm_x460_inr_Foreach.scala 74:112:@32126.4]
  wire [31:0] b454_number; // @[Math.scala 723:22:@32085.4 Math.scala 724:14:@32086.4]
  _ _ ( // @[Math.scala 720:24:@32080.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@32109.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@32118.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b455 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x460_inr_Foreach.scala 62:18:@32088.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x460_inr_Foreach.scala 67:129:@32092.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@32095.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x460_inr_Foreach.scala 67:146:@32096.4]
  assign x458_tuple = {1'h1,io_in_x243_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@32106.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32123.4 package.scala 96:25:@32124.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@32125.4]
  assign x579_b455_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@32114.4 package.scala 96:25:@32115.4]
  assign _T_293 = _T_292 & x579_b455_D2; // @[sm_x460_inr_Foreach.scala 74:112:@32126.4]
  assign b454_number = __io_result; // @[Math.scala 723:22:@32085.4 Math.scala 724:14:@32086.4]
  assign io_in_x243_outbuf_0_rPort_0_ofs_0 = b454_number[20:0]; // @[MemInterfaceType.scala 107:54:@32099.4]
  assign io_in_x243_outbuf_0_rPort_0_en_0 = _T_279 & b455; // @[MemInterfaceType.scala 110:79:@32101.4]
  assign io_in_x243_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32100.4]
  assign io_in_x445_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x460_inr_Foreach.scala 74:18:@32128.4]
  assign io_in_x445_bits_wdata_0 = x458_tuple[31:0]; // @[sm_x460_inr_Foreach.scala 75:26:@32130.4]
  assign io_in_x445_bits_wstrb = x458_tuple[32]; // @[sm_x460_inr_Foreach.scala 76:23:@32132.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@32083.4]
  assign RetimeWrapper_clock = clock; // @[:@32110.4]
  assign RetimeWrapper_reset = reset; // @[:@32111.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32113.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@32112.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32119.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32120.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32122.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32121.4]
endmodule
module x464_inr_UnitPipe_sm( // @[:@32288.2]
  input   clock, // @[:@32289.4]
  input   reset, // @[:@32290.4]
  input   io_enable, // @[:@32291.4]
  output  io_done, // @[:@32291.4]
  output  io_doneLatch, // @[:@32291.4]
  input   io_ctrDone, // @[:@32291.4]
  output  io_datapathEn, // @[:@32291.4]
  output  io_ctrInc, // @[:@32291.4]
  input   io_parentAck // @[:@32291.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@32293.4]
  wire  active_reset; // @[Controllers.scala 261:22:@32293.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@32293.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@32293.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@32293.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@32293.4]
  wire  done_clock; // @[Controllers.scala 262:20:@32296.4]
  wire  done_reset; // @[Controllers.scala 262:20:@32296.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@32296.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@32296.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@32296.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@32296.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32330.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32330.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32330.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32330.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32330.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32352.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32352.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32352.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32352.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32352.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32364.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32364.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32364.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32364.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32364.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32372.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32372.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32372.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32372.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32372.4]
  wire  _T_80; // @[Controllers.scala 264:48:@32301.4]
  wire  _T_81; // @[Controllers.scala 264:46:@32302.4]
  wire  _T_82; // @[Controllers.scala 264:62:@32303.4]
  wire  _T_100; // @[package.scala 100:49:@32321.4]
  reg  _T_103; // @[package.scala 48:56:@32322.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@32345.4]
  wire  _T_124; // @[package.scala 96:25:@32357.4 package.scala 96:25:@32358.4]
  wire  _T_126; // @[package.scala 100:49:@32359.4]
  reg  _T_129; // @[package.scala 48:56:@32360.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@32382.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@32384.4]
  reg  _T_153; // @[package.scala 48:56:@32385.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@32387.4]
  wire  _T_156; // @[Controllers.scala 292:61:@32388.4]
  wire  _T_157; // @[Controllers.scala 292:24:@32389.4]
  SRFF active ( // @[Controllers.scala 261:22:@32293.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@32296.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32330.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32352.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32364.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32372.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@32301.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@32302.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@32303.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@32321.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@32345.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32357.4 package.scala 96:25:@32358.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@32359.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@32384.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@32387.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@32388.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@32389.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@32363.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@32391.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@32348.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@32351.4]
  assign active_clock = clock; // @[:@32294.4]
  assign active_reset = reset; // @[:@32295.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@32306.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@32310.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@32311.4]
  assign done_clock = clock; // @[:@32297.4]
  assign done_reset = reset; // @[:@32298.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@32326.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@32319.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@32320.4]
  assign RetimeWrapper_clock = clock; // @[:@32331.4]
  assign RetimeWrapper_reset = reset; // @[:@32332.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32334.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@32333.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32353.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32354.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32356.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@32355.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32365.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32366.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32368.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@32367.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32373.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32374.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32376.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@32375.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1( // @[:@32466.2]
  output  io_in_x446_ready, // @[:@32469.4]
  input   io_sigsIn_datapathEn // @[:@32469.4]
);
  assign io_in_x446_ready = io_sigsIn_datapathEn; // @[sm_x464_inr_UnitPipe.scala 57:18:@32481.4]
endmodule
module x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1( // @[:@32484.2]
  input         clock, // @[:@32485.4]
  input         reset, // @[:@32486.4]
  output [20:0] io_in_x243_outbuf_0_rPort_0_ofs_0, // @[:@32487.4]
  output        io_in_x243_outbuf_0_rPort_0_en_0, // @[:@32487.4]
  output        io_in_x243_outbuf_0_rPort_0_backpressure, // @[:@32487.4]
  input  [31:0] io_in_x243_outbuf_0_rPort_0_output_0, // @[:@32487.4]
  input         io_in_x444_ready, // @[:@32487.4]
  output        io_in_x444_valid, // @[:@32487.4]
  output [63:0] io_in_x444_bits_addr, // @[:@32487.4]
  output [31:0] io_in_x444_bits_size, // @[:@32487.4]
  input         io_in_x445_ready, // @[:@32487.4]
  output        io_in_x445_valid, // @[:@32487.4]
  output [31:0] io_in_x445_bits_wdata_0, // @[:@32487.4]
  output        io_in_x445_bits_wstrb, // @[:@32487.4]
  output        io_in_x446_ready, // @[:@32487.4]
  input         io_in_x446_valid, // @[:@32487.4]
  input  [63:0] io_in_x239_outdram_number, // @[:@32487.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@32487.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@32487.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@32487.4]
  input         io_sigsIn_smChildAcks_0, // @[:@32487.4]
  input         io_sigsIn_smChildAcks_1, // @[:@32487.4]
  input         io_sigsIn_smChildAcks_2, // @[:@32487.4]
  output        io_sigsOut_smDoneIn_0, // @[:@32487.4]
  output        io_sigsOut_smDoneIn_1, // @[:@32487.4]
  output        io_sigsOut_smDoneIn_2, // @[:@32487.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@32487.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@32487.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@32487.4]
  input         io_rr // @[:@32487.4]
);
  wire  x451_inr_UnitPipe_sm_clock; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_reset; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_enable; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_done; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_doneLatch; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_ctrDone; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_datapathEn; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_ctrInc; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_parentAck; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  x451_inr_UnitPipe_sm_io_backpressure; // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32611.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32611.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32611.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32611.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32611.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32619.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32619.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32619.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32619.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32619.4]
  wire  x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_valid; // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
  wire [63:0] x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_bits_addr; // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
  wire [31:0] x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_bits_size; // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
  wire [63:0] x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x239_outdram_number; // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
  wire  x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
  wire  x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
  wire  x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_rr; // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
  wire  x453_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@32717.4]
  wire  x453_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@32717.4]
  wire  x453_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@32717.4]
  wire  x453_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@32717.4]
  wire [22:0] x453_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@32717.4]
  wire  x453_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@32717.4]
  wire  x453_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@32717.4]
  wire  x460_inr_Foreach_sm_clock; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_reset; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_enable; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_done; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_doneLatch; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_ctrDone; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_datapathEn; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_ctrInc; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_ctrRst; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_parentAck; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_backpressure; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  x460_inr_Foreach_sm_io_break; // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32798.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32798.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32798.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32798.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32798.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32838.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32838.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32838.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32838.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32838.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@32846.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@32846.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@32846.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@32846.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@32846.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_clock; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_reset; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire [20:0] x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_en_0; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire [31:0] x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_output_0; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_valid; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire [31:0] x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_bits_wdata_0; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_bits_wstrb; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire [31:0] x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_rr; // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
  wire  x464_inr_UnitPipe_sm_clock; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_reset; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_io_enable; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_io_done; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_io_doneLatch; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_io_ctrDone; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_io_datapathEn; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_io_ctrInc; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  x464_inr_UnitPipe_sm_io_parentAck; // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@33058.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@33066.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@33066.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@33066.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@33066.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@33066.4]
  wire  x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1_io_in_x446_ready; // @[sm_x464_inr_UnitPipe.scala 60:24:@33096.4]
  wire  x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x464_inr_UnitPipe.scala 60:24:@33096.4]
  wire  _T_359; // @[package.scala 100:49:@32582.4]
  reg  _T_362; // @[package.scala 48:56:@32583.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@32616.4 package.scala 96:25:@32617.4]
  wire  _T_381; // @[package.scala 96:25:@32624.4 package.scala 96:25:@32625.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@32627.4]
  wire  _T_454; // @[package.scala 96:25:@32803.4 package.scala 96:25:@32804.4]
  wire  _T_468; // @[package.scala 96:25:@32843.4 package.scala 96:25:@32844.4]
  wire  _T_474; // @[package.scala 96:25:@32851.4 package.scala 96:25:@32852.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@32854.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@32863.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@32864.4]
  wire  _T_547; // @[package.scala 100:49:@33029.4]
  reg  _T_550; // @[package.scala 48:56:@33030.4]
  reg [31:0] _RAND_1;
  wire  x464_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x465_outr_UnitPipe.scala 101:55:@33036.4]
  wire  _T_563; // @[package.scala 96:25:@33063.4 package.scala 96:25:@33064.4]
  wire  _T_569; // @[package.scala 96:25:@33071.4 package.scala 96:25:@33072.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@33074.4]
  wire  x464_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@33075.4]
  x451_inr_UnitPipe_sm x451_inr_UnitPipe_sm ( // @[sm_x451_inr_UnitPipe.scala 33:18:@32554.4]
    .clock(x451_inr_UnitPipe_sm_clock),
    .reset(x451_inr_UnitPipe_sm_reset),
    .io_enable(x451_inr_UnitPipe_sm_io_enable),
    .io_done(x451_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x451_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x451_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x451_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x451_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x451_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x451_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32611.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32619.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1 x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1 ( // @[sm_x451_inr_UnitPipe.scala 69:24:@32649.4]
    .io_in_x444_valid(x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_valid),
    .io_in_x444_bits_addr(x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_bits_addr),
    .io_in_x444_bits_size(x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_bits_size),
    .io_in_x239_outdram_number(x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x239_outdram_number),
    .io_sigsIn_backpressure(x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_rr)
  );
  x453_ctrchain x453_ctrchain ( // @[SpatialBlocks.scala 37:22:@32717.4]
    .clock(x453_ctrchain_clock),
    .reset(x453_ctrchain_reset),
    .io_input_reset(x453_ctrchain_io_input_reset),
    .io_input_enable(x453_ctrchain_io_input_enable),
    .io_output_counts_0(x453_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x453_ctrchain_io_output_oobs_0),
    .io_output_done(x453_ctrchain_io_output_done)
  );
  x460_inr_Foreach_sm x460_inr_Foreach_sm ( // @[sm_x460_inr_Foreach.scala 33:18:@32770.4]
    .clock(x460_inr_Foreach_sm_clock),
    .reset(x460_inr_Foreach_sm_reset),
    .io_enable(x460_inr_Foreach_sm_io_enable),
    .io_done(x460_inr_Foreach_sm_io_done),
    .io_doneLatch(x460_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x460_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x460_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x460_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x460_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x460_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x460_inr_Foreach_sm_io_backpressure),
    .io_break(x460_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32798.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32838.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@32846.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x460_inr_Foreach_kernelx460_inr_Foreach_concrete1 x460_inr_Foreach_kernelx460_inr_Foreach_concrete1 ( // @[sm_x460_inr_Foreach.scala 78:24:@32881.4]
    .clock(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_clock),
    .reset(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_reset),
    .io_in_x243_outbuf_0_rPort_0_ofs_0(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0),
    .io_in_x243_outbuf_0_rPort_0_en_0(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_en_0),
    .io_in_x243_outbuf_0_rPort_0_backpressure(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure),
    .io_in_x243_outbuf_0_rPort_0_output_0(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_output_0),
    .io_in_x445_valid(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_valid),
    .io_in_x445_bits_wdata_0(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_bits_wdata_0),
    .io_in_x445_bits_wstrb(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_bits_wstrb),
    .io_sigsIn_backpressure(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_rr)
  );
  x464_inr_UnitPipe_sm x464_inr_UnitPipe_sm ( // @[sm_x464_inr_UnitPipe.scala 32:18:@33001.4]
    .clock(x464_inr_UnitPipe_sm_clock),
    .reset(x464_inr_UnitPipe_sm_reset),
    .io_enable(x464_inr_UnitPipe_sm_io_enable),
    .io_done(x464_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x464_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x464_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x464_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x464_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x464_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@33058.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@33066.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1 x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1 ( // @[sm_x464_inr_UnitPipe.scala 60:24:@33096.4]
    .io_in_x446_ready(x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1_io_in_x446_ready),
    .io_sigsIn_datapathEn(x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x451_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@32582.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@32616.4 package.scala 96:25:@32617.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32624.4 package.scala 96:25:@32625.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@32627.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@32803.4 package.scala 96:25:@32804.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@32843.4 package.scala 96:25:@32844.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@32851.4 package.scala 96:25:@32852.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@32854.4]
  assign _T_479 = x460_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@32863.4]
  assign _T_480 = ~ x460_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@32864.4]
  assign _T_547 = x464_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33029.4]
  assign x464_inr_UnitPipe_sigsIn_forwardpressure = io_in_x446_valid | x464_inr_UnitPipe_sm_io_doneLatch; // @[sm_x465_outr_UnitPipe.scala 101:55:@33036.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@33063.4 package.scala 96:25:@33064.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@33071.4 package.scala 96:25:@33072.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@33074.4]
  assign x464_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@33075.4]
  assign io_in_x243_outbuf_0_rPort_0_ofs_0 = x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@32932.4]
  assign io_in_x243_outbuf_0_rPort_0_en_0 = x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@32931.4]
  assign io_in_x243_outbuf_0_rPort_0_backpressure = x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@32930.4]
  assign io_in_x444_valid = x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_valid; // @[sm_x451_inr_UnitPipe.scala 49:23:@32687.4]
  assign io_in_x444_bits_addr = x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_bits_addr; // @[sm_x451_inr_UnitPipe.scala 49:23:@32686.4]
  assign io_in_x444_bits_size = x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x444_bits_size; // @[sm_x451_inr_UnitPipe.scala 49:23:@32685.4]
  assign io_in_x445_valid = x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_valid; // @[sm_x460_inr_Foreach.scala 50:23:@32936.4]
  assign io_in_x445_bits_wdata_0 = x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_bits_wdata_0; // @[sm_x460_inr_Foreach.scala 50:23:@32935.4]
  assign io_in_x445_bits_wstrb = x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x445_bits_wstrb; // @[sm_x460_inr_Foreach.scala 50:23:@32934.4]
  assign io_in_x446_ready = x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1_io_in_x446_ready; // @[sm_x464_inr_UnitPipe.scala 46:23:@33132.4]
  assign io_sigsOut_smDoneIn_0 = x451_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@32634.4]
  assign io_sigsOut_smDoneIn_1 = x460_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@32861.4]
  assign io_sigsOut_smDoneIn_2 = x464_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33081.4]
  assign io_sigsOut_smCtrCopyDone_0 = x451_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@32648.4]
  assign io_sigsOut_smCtrCopyDone_1 = x460_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@32880.4]
  assign io_sigsOut_smCtrCopyDone_2 = x464_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@33095.4]
  assign x451_inr_UnitPipe_sm_clock = clock; // @[:@32555.4]
  assign x451_inr_UnitPipe_sm_reset = reset; // @[:@32556.4]
  assign x451_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@32631.4]
  assign x451_inr_UnitPipe_sm_io_ctrDone = x451_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x465_outr_UnitPipe.scala 77:39:@32586.4]
  assign x451_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@32633.4]
  assign x451_inr_UnitPipe_sm_io_backpressure = io_in_x444_ready | x451_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@32605.4]
  assign RetimeWrapper_clock = clock; // @[:@32612.4]
  assign RetimeWrapper_reset = reset; // @[:@32613.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32615.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@32614.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32620.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32621.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32623.4]
  assign RetimeWrapper_1_io_in = x451_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@32622.4]
  assign x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_in_x239_outdram_number = io_in_x239_outdram_number; // @[sm_x451_inr_UnitPipe.scala 50:31:@32689.4]
  assign x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x444_ready | x451_inr_UnitPipe_sm_io_doneLatch; // @[sm_x451_inr_UnitPipe.scala 74:22:@32704.4]
  assign x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x451_inr_UnitPipe_sm_io_datapathEn; // @[sm_x451_inr_UnitPipe.scala 74:22:@32702.4]
  assign x451_inr_UnitPipe_kernelx451_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x451_inr_UnitPipe.scala 73:18:@32690.4]
  assign x453_ctrchain_clock = clock; // @[:@32718.4]
  assign x453_ctrchain_reset = reset; // @[:@32719.4]
  assign x453_ctrchain_io_input_reset = x460_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@32879.4]
  assign x453_ctrchain_io_input_enable = x460_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@32831.4 SpatialBlocks.scala 159:42:@32878.4]
  assign x460_inr_Foreach_sm_clock = clock; // @[:@32771.4]
  assign x460_inr_Foreach_sm_reset = reset; // @[:@32772.4]
  assign x460_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@32858.4]
  assign x460_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x465_outr_UnitPipe.scala 90:38:@32806.4]
  assign x460_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@32860.4]
  assign x460_inr_Foreach_sm_io_backpressure = io_in_x445_ready | x460_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@32832.4]
  assign x460_inr_Foreach_sm_io_break = 1'h0; // @[sm_x465_outr_UnitPipe.scala 94:36:@32812.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32799.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32800.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32802.4]
  assign RetimeWrapper_2_io_in = x453_ctrchain_io_output_done; // @[package.scala 94:16:@32801.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32839.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32840.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32842.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@32841.4]
  assign RetimeWrapper_4_clock = clock; // @[:@32847.4]
  assign RetimeWrapper_4_reset = reset; // @[:@32848.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@32850.4]
  assign RetimeWrapper_4_io_in = x460_inr_Foreach_sm_io_done; // @[package.scala 94:16:@32849.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_clock = clock; // @[:@32882.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_reset = reset; // @[:@32883.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_in_x243_outbuf_0_rPort_0_output_0 = io_in_x243_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@32929.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x445_ready | x460_inr_Foreach_sm_io_doneLatch; // @[sm_x460_inr_Foreach.scala 83:22:@32952.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x460_inr_Foreach.scala 83:22:@32950.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_break = x460_inr_Foreach_sm_io_break; // @[sm_x460_inr_Foreach.scala 83:22:@32948.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x453_ctrchain_io_output_counts_0[22]}},x453_ctrchain_io_output_counts_0}; // @[sm_x460_inr_Foreach.scala 83:22:@32943.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x453_ctrchain_io_output_oobs_0; // @[sm_x460_inr_Foreach.scala 83:22:@32942.4]
  assign x460_inr_Foreach_kernelx460_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x460_inr_Foreach.scala 82:18:@32938.4]
  assign x464_inr_UnitPipe_sm_clock = clock; // @[:@33002.4]
  assign x464_inr_UnitPipe_sm_reset = reset; // @[:@33003.4]
  assign x464_inr_UnitPipe_sm_io_enable = x464_inr_UnitPipe_sigsIn_baseEn & x464_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@33078.4]
  assign x464_inr_UnitPipe_sm_io_ctrDone = x464_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x465_outr_UnitPipe.scala 99:39:@33033.4]
  assign x464_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@33080.4]
  assign RetimeWrapper_5_clock = clock; // @[:@33059.4]
  assign RetimeWrapper_5_reset = reset; // @[:@33060.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@33062.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@33061.4]
  assign RetimeWrapper_6_clock = clock; // @[:@33067.4]
  assign RetimeWrapper_6_reset = reset; // @[:@33068.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@33070.4]
  assign RetimeWrapper_6_io_in = x464_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33069.4]
  assign x464_inr_UnitPipe_kernelx464_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x464_inr_UnitPipe_sm_io_datapathEn; // @[sm_x464_inr_UnitPipe.scala 65:22:@33145.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x518_kernelx518_concrete1( // @[:@33161.2]
  input          clock, // @[:@33162.4]
  input          reset, // @[:@33163.4]
  output [20:0]  io_in_x243_outbuf_0_rPort_0_ofs_0, // @[:@33164.4]
  output         io_in_x243_outbuf_0_rPort_0_en_0, // @[:@33164.4]
  output         io_in_x243_outbuf_0_rPort_0_backpressure, // @[:@33164.4]
  input  [31:0]  io_in_x243_outbuf_0_rPort_0_output_0, // @[:@33164.4]
  input          io_in_x444_ready, // @[:@33164.4]
  output         io_in_x444_valid, // @[:@33164.4]
  output [63:0]  io_in_x444_bits_addr, // @[:@33164.4]
  output [31:0]  io_in_x444_bits_size, // @[:@33164.4]
  input          io_in_x445_ready, // @[:@33164.4]
  output         io_in_x445_valid, // @[:@33164.4]
  output [31:0]  io_in_x445_bits_wdata_0, // @[:@33164.4]
  output         io_in_x445_bits_wstrb, // @[:@33164.4]
  input          io_in_x241_TVALID, // @[:@33164.4]
  output         io_in_x241_TREADY, // @[:@33164.4]
  input  [255:0] io_in_x241_TDATA, // @[:@33164.4]
  input  [7:0]   io_in_x241_TID, // @[:@33164.4]
  input  [7:0]   io_in_x241_TDEST, // @[:@33164.4]
  output         io_in_x446_ready, // @[:@33164.4]
  input          io_in_x446_valid, // @[:@33164.4]
  input  [63:0]  io_in_x239_outdram_number, // @[:@33164.4]
  output         io_in_x242_TVALID, // @[:@33164.4]
  input          io_in_x242_TREADY, // @[:@33164.4]
  output [255:0] io_in_x242_TDATA, // @[:@33164.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@33164.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@33164.4]
  input          io_sigsIn_smChildAcks_0, // @[:@33164.4]
  input          io_sigsIn_smChildAcks_1, // @[:@33164.4]
  output         io_sigsOut_smDoneIn_0, // @[:@33164.4]
  output         io_sigsOut_smDoneIn_1, // @[:@33164.4]
  input          io_rr // @[:@33164.4]
);
  wire  x443_outr_UnitPipe_sm_clock; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_reset; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_enable; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_done; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_parentAck; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_childAck_0; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_childAck_1; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  x443_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33299.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33299.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33299.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33299.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33299.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33307.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33307.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33307.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33307.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33307.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_clock; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_reset; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TVALID; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TREADY; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire [255:0] x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TDATA; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire [7:0] x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TID; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire [7:0] x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TDEST; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TVALID; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TREADY; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire [255:0] x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TDATA; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_rr; // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
  wire  x465_outr_UnitPipe_sm_clock; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_reset; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_enable; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_done; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_parentAck; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_childAck_0; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_childAck_1; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_childAck_2; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  x465_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@33588.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@33588.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@33588.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@33588.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@33588.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@33596.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@33596.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@33596.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@33596.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@33596.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_clock; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_reset; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire [20:0] x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_en_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire [31:0] x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_output_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_ready; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_valid; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire [63:0] x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_bits_addr; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire [31:0] x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_bits_size; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_ready; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_valid; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire [31:0] x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_bits_wdata_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_bits_wstrb; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x446_ready; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x446_valid; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire [63:0] x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x239_outdram_number; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_rr; // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
  wire  _T_408; // @[package.scala 96:25:@33304.4 package.scala 96:25:@33305.4]
  wire  _T_414; // @[package.scala 96:25:@33312.4 package.scala 96:25:@33313.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@33315.4]
  wire  _T_508; // @[package.scala 96:25:@33593.4 package.scala 96:25:@33594.4]
  wire  _T_514; // @[package.scala 96:25:@33601.4 package.scala 96:25:@33602.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@33604.4]
  x443_outr_UnitPipe_sm x443_outr_UnitPipe_sm ( // @[sm_x443_outr_UnitPipe.scala 32:18:@33237.4]
    .clock(x443_outr_UnitPipe_sm_clock),
    .reset(x443_outr_UnitPipe_sm_reset),
    .io_enable(x443_outr_UnitPipe_sm_io_enable),
    .io_done(x443_outr_UnitPipe_sm_io_done),
    .io_parentAck(x443_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x443_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x443_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x443_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x443_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x443_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x443_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x443_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x443_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33299.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33307.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1 x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1 ( // @[sm_x443_outr_UnitPipe.scala 87:24:@33338.4]
    .clock(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_clock),
    .reset(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_reset),
    .io_in_x241_TVALID(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TVALID),
    .io_in_x241_TREADY(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TREADY),
    .io_in_x241_TDATA(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TDATA),
    .io_in_x241_TID(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TID),
    .io_in_x241_TDEST(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TDEST),
    .io_in_x242_TVALID(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TVALID),
    .io_in_x242_TREADY(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TREADY),
    .io_in_x242_TDATA(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TDATA),
    .io_sigsIn_smEnableOuts_0(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_rr)
  );
  x465_outr_UnitPipe_sm x465_outr_UnitPipe_sm ( // @[sm_x465_outr_UnitPipe.scala 36:18:@33516.4]
    .clock(x465_outr_UnitPipe_sm_clock),
    .reset(x465_outr_UnitPipe_sm_reset),
    .io_enable(x465_outr_UnitPipe_sm_io_enable),
    .io_done(x465_outr_UnitPipe_sm_io_done),
    .io_parentAck(x465_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x465_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x465_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x465_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x465_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x465_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x465_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x465_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x465_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x465_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x465_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x465_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x465_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@33588.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@33596.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1 x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1 ( // @[sm_x465_outr_UnitPipe.scala 108:24:@33628.4]
    .clock(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_clock),
    .reset(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_reset),
    .io_in_x243_outbuf_0_rPort_0_ofs_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0),
    .io_in_x243_outbuf_0_rPort_0_en_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_en_0),
    .io_in_x243_outbuf_0_rPort_0_backpressure(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure),
    .io_in_x243_outbuf_0_rPort_0_output_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_output_0),
    .io_in_x444_ready(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_ready),
    .io_in_x444_valid(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_valid),
    .io_in_x444_bits_addr(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_bits_addr),
    .io_in_x444_bits_size(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_bits_size),
    .io_in_x445_ready(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_ready),
    .io_in_x445_valid(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_valid),
    .io_in_x445_bits_wdata_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_bits_wdata_0),
    .io_in_x445_bits_wstrb(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_bits_wstrb),
    .io_in_x446_ready(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x446_ready),
    .io_in_x446_valid(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x446_valid),
    .io_in_x239_outdram_number(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x239_outdram_number),
    .io_sigsIn_smEnableOuts_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@33304.4 package.scala 96:25:@33305.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33312.4 package.scala 96:25:@33313.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@33315.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@33593.4 package.scala 96:25:@33594.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@33601.4 package.scala 96:25:@33602.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@33604.4]
  assign io_in_x243_outbuf_0_rPort_0_ofs_0 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@33711.4]
  assign io_in_x243_outbuf_0_rPort_0_en_0 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@33710.4]
  assign io_in_x243_outbuf_0_rPort_0_backpressure = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@33709.4]
  assign io_in_x444_valid = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_valid; // @[sm_x465_outr_UnitPipe.scala 59:23:@33715.4]
  assign io_in_x444_bits_addr = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_bits_addr; // @[sm_x465_outr_UnitPipe.scala 59:23:@33714.4]
  assign io_in_x444_bits_size = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_bits_size; // @[sm_x465_outr_UnitPipe.scala 59:23:@33713.4]
  assign io_in_x445_valid = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_valid; // @[sm_x465_outr_UnitPipe.scala 60:23:@33719.4]
  assign io_in_x445_bits_wdata_0 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_bits_wdata_0; // @[sm_x465_outr_UnitPipe.scala 60:23:@33718.4]
  assign io_in_x445_bits_wstrb = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_bits_wstrb; // @[sm_x465_outr_UnitPipe.scala 60:23:@33717.4]
  assign io_in_x241_TREADY = x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TREADY; // @[sm_x443_outr_UnitPipe.scala 48:23:@33406.4]
  assign io_in_x446_ready = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x446_ready; // @[sm_x465_outr_UnitPipe.scala 61:23:@33723.4]
  assign io_in_x242_TVALID = x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TVALID; // @[sm_x443_outr_UnitPipe.scala 49:23:@33416.4]
  assign io_in_x242_TDATA = x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TDATA; // @[sm_x443_outr_UnitPipe.scala 49:23:@33414.4]
  assign io_sigsOut_smDoneIn_0 = x443_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33322.4]
  assign io_sigsOut_smDoneIn_1 = x465_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33611.4]
  assign x443_outr_UnitPipe_sm_clock = clock; // @[:@33238.4]
  assign x443_outr_UnitPipe_sm_reset = reset; // @[:@33239.4]
  assign x443_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@33319.4]
  assign x443_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@33321.4]
  assign x443_outr_UnitPipe_sm_io_doneIn_0 = x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33289.4]
  assign x443_outr_UnitPipe_sm_io_doneIn_1 = x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33290.4]
  assign x443_outr_UnitPipe_sm_io_ctrCopyDone_0 = x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@33336.4]
  assign x443_outr_UnitPipe_sm_io_ctrCopyDone_1 = x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@33337.4]
  assign RetimeWrapper_clock = clock; // @[:@33300.4]
  assign RetimeWrapper_reset = reset; // @[:@33301.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33303.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@33302.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33308.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33309.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33311.4]
  assign RetimeWrapper_1_io_in = x443_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33310.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_clock = clock; // @[:@33339.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_reset = reset; // @[:@33340.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TVALID = io_in_x241_TVALID; // @[sm_x443_outr_UnitPipe.scala 48:23:@33407.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TDATA = io_in_x241_TDATA; // @[sm_x443_outr_UnitPipe.scala 48:23:@33405.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TID = io_in_x241_TID; // @[sm_x443_outr_UnitPipe.scala 48:23:@33401.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x241_TDEST = io_in_x241_TDEST; // @[sm_x443_outr_UnitPipe.scala 48:23:@33400.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_in_x242_TREADY = io_in_x242_TREADY; // @[sm_x443_outr_UnitPipe.scala 49:23:@33415.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x443_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x443_outr_UnitPipe.scala 92:22:@33432.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x443_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x443_outr_UnitPipe.scala 92:22:@33433.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x443_outr_UnitPipe_sm_io_childAck_0; // @[sm_x443_outr_UnitPipe.scala 92:22:@33428.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x443_outr_UnitPipe_sm_io_childAck_1; // @[sm_x443_outr_UnitPipe.scala 92:22:@33429.4]
  assign x443_outr_UnitPipe_kernelx443_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x443_outr_UnitPipe.scala 91:18:@33417.4]
  assign x465_outr_UnitPipe_sm_clock = clock; // @[:@33517.4]
  assign x465_outr_UnitPipe_sm_reset = reset; // @[:@33518.4]
  assign x465_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@33608.4]
  assign x465_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@33610.4]
  assign x465_outr_UnitPipe_sm_io_doneIn_0 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33576.4]
  assign x465_outr_UnitPipe_sm_io_doneIn_1 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33577.4]
  assign x465_outr_UnitPipe_sm_io_doneIn_2 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@33578.4]
  assign x465_outr_UnitPipe_sm_io_ctrCopyDone_0 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@33625.4]
  assign x465_outr_UnitPipe_sm_io_ctrCopyDone_1 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@33626.4]
  assign x465_outr_UnitPipe_sm_io_ctrCopyDone_2 = x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@33627.4]
  assign RetimeWrapper_2_clock = clock; // @[:@33589.4]
  assign RetimeWrapper_2_reset = reset; // @[:@33590.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@33592.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@33591.4]
  assign RetimeWrapper_3_clock = clock; // @[:@33597.4]
  assign RetimeWrapper_3_reset = reset; // @[:@33598.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@33600.4]
  assign RetimeWrapper_3_io_in = x465_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33599.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_clock = clock; // @[:@33629.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_reset = reset; // @[:@33630.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x243_outbuf_0_rPort_0_output_0 = io_in_x243_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@33708.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x444_ready = io_in_x444_ready; // @[sm_x465_outr_UnitPipe.scala 59:23:@33716.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x445_ready = io_in_x445_ready; // @[sm_x465_outr_UnitPipe.scala 60:23:@33720.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x446_valid = io_in_x446_valid; // @[sm_x465_outr_UnitPipe.scala 61:23:@33722.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_in_x239_outdram_number = io_in_x239_outdram_number; // @[sm_x465_outr_UnitPipe.scala 62:31:@33724.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x465_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x465_outr_UnitPipe.scala 113:22:@33747.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x465_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x465_outr_UnitPipe.scala 113:22:@33748.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x465_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x465_outr_UnitPipe.scala 113:22:@33749.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x465_outr_UnitPipe_sm_io_childAck_0; // @[sm_x465_outr_UnitPipe.scala 113:22:@33741.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x465_outr_UnitPipe_sm_io_childAck_1; // @[sm_x465_outr_UnitPipe.scala 113:22:@33742.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x465_outr_UnitPipe_sm_io_childAck_2; // @[sm_x465_outr_UnitPipe.scala 113:22:@33743.4]
  assign x465_outr_UnitPipe_kernelx465_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x465_outr_UnitPipe.scala 112:18:@33725.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@33777.2]
  input          clock, // @[:@33778.4]
  input          reset, // @[:@33779.4]
  input          io_in_x444_ready, // @[:@33780.4]
  output         io_in_x444_valid, // @[:@33780.4]
  output [63:0]  io_in_x444_bits_addr, // @[:@33780.4]
  output [31:0]  io_in_x444_bits_size, // @[:@33780.4]
  input          io_in_x445_ready, // @[:@33780.4]
  output         io_in_x445_valid, // @[:@33780.4]
  output [31:0]  io_in_x445_bits_wdata_0, // @[:@33780.4]
  output         io_in_x445_bits_wstrb, // @[:@33780.4]
  input          io_in_x241_TVALID, // @[:@33780.4]
  output         io_in_x241_TREADY, // @[:@33780.4]
  input  [255:0] io_in_x241_TDATA, // @[:@33780.4]
  input  [7:0]   io_in_x241_TID, // @[:@33780.4]
  input  [7:0]   io_in_x241_TDEST, // @[:@33780.4]
  output         io_in_x446_ready, // @[:@33780.4]
  input          io_in_x446_valid, // @[:@33780.4]
  input  [63:0]  io_in_x239_outdram_number, // @[:@33780.4]
  output         io_in_x242_TVALID, // @[:@33780.4]
  input          io_in_x242_TREADY, // @[:@33780.4]
  output [255:0] io_in_x242_TDATA, // @[:@33780.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@33780.4]
  input          io_sigsIn_smChildAcks_0, // @[:@33780.4]
  output         io_sigsOut_smDoneIn_0, // @[:@33780.4]
  input          io_rr // @[:@33780.4]
);
  wire  x243_outbuf_0_clock; // @[m_x243_outbuf_0.scala 27:17:@33790.4]
  wire  x243_outbuf_0_reset; // @[m_x243_outbuf_0.scala 27:17:@33790.4]
  wire [20:0] x243_outbuf_0_io_rPort_0_ofs_0; // @[m_x243_outbuf_0.scala 27:17:@33790.4]
  wire  x243_outbuf_0_io_rPort_0_en_0; // @[m_x243_outbuf_0.scala 27:17:@33790.4]
  wire  x243_outbuf_0_io_rPort_0_backpressure; // @[m_x243_outbuf_0.scala 27:17:@33790.4]
  wire [31:0] x243_outbuf_0_io_rPort_0_output_0; // @[m_x243_outbuf_0.scala 27:17:@33790.4]
  wire  x518_sm_clock; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_reset; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_enable; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_done; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_ctrDone; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_ctrInc; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_parentAck; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_doneIn_0; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_doneIn_1; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_enableOut_0; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_enableOut_1; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_childAck_0; // @[sm_x518.scala 37:18:@33848.4]
  wire  x518_sm_io_childAck_1; // @[sm_x518.scala 37:18:@33848.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33915.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33915.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33915.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33915.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33915.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33923.4]
  wire  x518_kernelx518_concrete1_clock; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_reset; // @[sm_x518.scala 102:24:@33952.4]
  wire [20:0] x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_en_0; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure; // @[sm_x518.scala 102:24:@33952.4]
  wire [31:0] x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_output_0; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x444_ready; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x444_valid; // @[sm_x518.scala 102:24:@33952.4]
  wire [63:0] x518_kernelx518_concrete1_io_in_x444_bits_addr; // @[sm_x518.scala 102:24:@33952.4]
  wire [31:0] x518_kernelx518_concrete1_io_in_x444_bits_size; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x445_ready; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x445_valid; // @[sm_x518.scala 102:24:@33952.4]
  wire [31:0] x518_kernelx518_concrete1_io_in_x445_bits_wdata_0; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x445_bits_wstrb; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x241_TVALID; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x241_TREADY; // @[sm_x518.scala 102:24:@33952.4]
  wire [255:0] x518_kernelx518_concrete1_io_in_x241_TDATA; // @[sm_x518.scala 102:24:@33952.4]
  wire [7:0] x518_kernelx518_concrete1_io_in_x241_TID; // @[sm_x518.scala 102:24:@33952.4]
  wire [7:0] x518_kernelx518_concrete1_io_in_x241_TDEST; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x446_ready; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x446_valid; // @[sm_x518.scala 102:24:@33952.4]
  wire [63:0] x518_kernelx518_concrete1_io_in_x239_outdram_number; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x242_TVALID; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_in_x242_TREADY; // @[sm_x518.scala 102:24:@33952.4]
  wire [255:0] x518_kernelx518_concrete1_io_in_x242_TDATA; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x518.scala 102:24:@33952.4]
  wire  x518_kernelx518_concrete1_io_rr; // @[sm_x518.scala 102:24:@33952.4]
  wire  _T_266; // @[package.scala 100:49:@33881.4]
  reg  _T_269; // @[package.scala 48:56:@33882.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@33920.4 package.scala 96:25:@33921.4]
  wire  _T_289; // @[package.scala 96:25:@33928.4 package.scala 96:25:@33929.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@33931.4]
  x243_outbuf_0 x243_outbuf_0 ( // @[m_x243_outbuf_0.scala 27:17:@33790.4]
    .clock(x243_outbuf_0_clock),
    .reset(x243_outbuf_0_reset),
    .io_rPort_0_ofs_0(x243_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x243_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x243_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x243_outbuf_0_io_rPort_0_output_0)
  );
  x518_sm x518_sm ( // @[sm_x518.scala 37:18:@33848.4]
    .clock(x518_sm_clock),
    .reset(x518_sm_reset),
    .io_enable(x518_sm_io_enable),
    .io_done(x518_sm_io_done),
    .io_ctrDone(x518_sm_io_ctrDone),
    .io_ctrInc(x518_sm_io_ctrInc),
    .io_parentAck(x518_sm_io_parentAck),
    .io_doneIn_0(x518_sm_io_doneIn_0),
    .io_doneIn_1(x518_sm_io_doneIn_1),
    .io_enableOut_0(x518_sm_io_enableOut_0),
    .io_enableOut_1(x518_sm_io_enableOut_1),
    .io_childAck_0(x518_sm_io_childAck_0),
    .io_childAck_1(x518_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33915.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33923.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x518_kernelx518_concrete1 x518_kernelx518_concrete1 ( // @[sm_x518.scala 102:24:@33952.4]
    .clock(x518_kernelx518_concrete1_clock),
    .reset(x518_kernelx518_concrete1_reset),
    .io_in_x243_outbuf_0_rPort_0_ofs_0(x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0),
    .io_in_x243_outbuf_0_rPort_0_en_0(x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_en_0),
    .io_in_x243_outbuf_0_rPort_0_backpressure(x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure),
    .io_in_x243_outbuf_0_rPort_0_output_0(x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_output_0),
    .io_in_x444_ready(x518_kernelx518_concrete1_io_in_x444_ready),
    .io_in_x444_valid(x518_kernelx518_concrete1_io_in_x444_valid),
    .io_in_x444_bits_addr(x518_kernelx518_concrete1_io_in_x444_bits_addr),
    .io_in_x444_bits_size(x518_kernelx518_concrete1_io_in_x444_bits_size),
    .io_in_x445_ready(x518_kernelx518_concrete1_io_in_x445_ready),
    .io_in_x445_valid(x518_kernelx518_concrete1_io_in_x445_valid),
    .io_in_x445_bits_wdata_0(x518_kernelx518_concrete1_io_in_x445_bits_wdata_0),
    .io_in_x445_bits_wstrb(x518_kernelx518_concrete1_io_in_x445_bits_wstrb),
    .io_in_x241_TVALID(x518_kernelx518_concrete1_io_in_x241_TVALID),
    .io_in_x241_TREADY(x518_kernelx518_concrete1_io_in_x241_TREADY),
    .io_in_x241_TDATA(x518_kernelx518_concrete1_io_in_x241_TDATA),
    .io_in_x241_TID(x518_kernelx518_concrete1_io_in_x241_TID),
    .io_in_x241_TDEST(x518_kernelx518_concrete1_io_in_x241_TDEST),
    .io_in_x446_ready(x518_kernelx518_concrete1_io_in_x446_ready),
    .io_in_x446_valid(x518_kernelx518_concrete1_io_in_x446_valid),
    .io_in_x239_outdram_number(x518_kernelx518_concrete1_io_in_x239_outdram_number),
    .io_in_x242_TVALID(x518_kernelx518_concrete1_io_in_x242_TVALID),
    .io_in_x242_TREADY(x518_kernelx518_concrete1_io_in_x242_TREADY),
    .io_in_x242_TDATA(x518_kernelx518_concrete1_io_in_x242_TDATA),
    .io_sigsIn_smEnableOuts_0(x518_kernelx518_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x518_kernelx518_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x518_kernelx518_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x518_kernelx518_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x518_kernelx518_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x518_kernelx518_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x518_kernelx518_concrete1_io_rr)
  );
  assign _T_266 = x518_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33881.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@33920.4 package.scala 96:25:@33921.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33928.4 package.scala 96:25:@33929.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@33931.4]
  assign io_in_x444_valid = x518_kernelx518_concrete1_io_in_x444_valid; // @[sm_x518.scala 64:23:@34038.4]
  assign io_in_x444_bits_addr = x518_kernelx518_concrete1_io_in_x444_bits_addr; // @[sm_x518.scala 64:23:@34037.4]
  assign io_in_x444_bits_size = x518_kernelx518_concrete1_io_in_x444_bits_size; // @[sm_x518.scala 64:23:@34036.4]
  assign io_in_x445_valid = x518_kernelx518_concrete1_io_in_x445_valid; // @[sm_x518.scala 65:23:@34042.4]
  assign io_in_x445_bits_wdata_0 = x518_kernelx518_concrete1_io_in_x445_bits_wdata_0; // @[sm_x518.scala 65:23:@34041.4]
  assign io_in_x445_bits_wstrb = x518_kernelx518_concrete1_io_in_x445_bits_wstrb; // @[sm_x518.scala 65:23:@34040.4]
  assign io_in_x241_TREADY = x518_kernelx518_concrete1_io_in_x241_TREADY; // @[sm_x518.scala 66:23:@34051.4]
  assign io_in_x446_ready = x518_kernelx518_concrete1_io_in_x446_ready; // @[sm_x518.scala 67:23:@34055.4]
  assign io_in_x242_TVALID = x518_kernelx518_concrete1_io_in_x242_TVALID; // @[sm_x518.scala 69:23:@34065.4]
  assign io_in_x242_TDATA = x518_kernelx518_concrete1_io_in_x242_TDATA; // @[sm_x518.scala 69:23:@34063.4]
  assign io_sigsOut_smDoneIn_0 = x518_sm_io_done; // @[SpatialBlocks.scala 156:53:@33938.4]
  assign x243_outbuf_0_clock = clock; // @[:@33791.4]
  assign x243_outbuf_0_reset = reset; // @[:@33792.4]
  assign x243_outbuf_0_io_rPort_0_ofs_0 = x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@34034.4]
  assign x243_outbuf_0_io_rPort_0_en_0 = x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@34033.4]
  assign x243_outbuf_0_io_rPort_0_backpressure = x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@34032.4]
  assign x518_sm_clock = clock; // @[:@33849.4]
  assign x518_sm_reset = reset; // @[:@33850.4]
  assign x518_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@33935.4]
  assign x518_sm_io_ctrDone = x518_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@33885.4]
  assign x518_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@33937.4]
  assign x518_sm_io_doneIn_0 = x518_kernelx518_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33905.4]
  assign x518_sm_io_doneIn_1 = x518_kernelx518_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33906.4]
  assign RetimeWrapper_clock = clock; // @[:@33916.4]
  assign RetimeWrapper_reset = reset; // @[:@33917.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33919.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@33918.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33924.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33925.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33927.4]
  assign RetimeWrapper_1_io_in = x518_sm_io_done; // @[package.scala 94:16:@33926.4]
  assign x518_kernelx518_concrete1_clock = clock; // @[:@33953.4]
  assign x518_kernelx518_concrete1_reset = reset; // @[:@33954.4]
  assign x518_kernelx518_concrete1_io_in_x243_outbuf_0_rPort_0_output_0 = x243_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@34031.4]
  assign x518_kernelx518_concrete1_io_in_x444_ready = io_in_x444_ready; // @[sm_x518.scala 64:23:@34039.4]
  assign x518_kernelx518_concrete1_io_in_x445_ready = io_in_x445_ready; // @[sm_x518.scala 65:23:@34043.4]
  assign x518_kernelx518_concrete1_io_in_x241_TVALID = io_in_x241_TVALID; // @[sm_x518.scala 66:23:@34052.4]
  assign x518_kernelx518_concrete1_io_in_x241_TDATA = io_in_x241_TDATA; // @[sm_x518.scala 66:23:@34050.4]
  assign x518_kernelx518_concrete1_io_in_x241_TID = io_in_x241_TID; // @[sm_x518.scala 66:23:@34046.4]
  assign x518_kernelx518_concrete1_io_in_x241_TDEST = io_in_x241_TDEST; // @[sm_x518.scala 66:23:@34045.4]
  assign x518_kernelx518_concrete1_io_in_x446_valid = io_in_x446_valid; // @[sm_x518.scala 67:23:@34054.4]
  assign x518_kernelx518_concrete1_io_in_x239_outdram_number = io_in_x239_outdram_number; // @[sm_x518.scala 68:31:@34056.4]
  assign x518_kernelx518_concrete1_io_in_x242_TREADY = io_in_x242_TREADY; // @[sm_x518.scala 69:23:@34064.4]
  assign x518_kernelx518_concrete1_io_sigsIn_smEnableOuts_0 = x518_sm_io_enableOut_0; // @[sm_x518.scala 107:22:@34076.4]
  assign x518_kernelx518_concrete1_io_sigsIn_smEnableOuts_1 = x518_sm_io_enableOut_1; // @[sm_x518.scala 107:22:@34077.4]
  assign x518_kernelx518_concrete1_io_sigsIn_smChildAcks_0 = x518_sm_io_childAck_0; // @[sm_x518.scala 107:22:@34072.4]
  assign x518_kernelx518_concrete1_io_sigsIn_smChildAcks_1 = x518_sm_io_childAck_1; // @[sm_x518.scala 107:22:@34073.4]
  assign x518_kernelx518_concrete1_io_rr = io_rr; // @[sm_x518.scala 106:18:@34066.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@34099.2]
  input          clock, // @[:@34100.4]
  input          reset, // @[:@34101.4]
  input          io_enable, // @[:@34102.4]
  output         io_done, // @[:@34102.4]
  input          io_reset, // @[:@34102.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@34102.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@34102.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@34102.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@34102.4]
  output         io_memStreams_loads_0_data_ready, // @[:@34102.4]
  input          io_memStreams_loads_0_data_valid, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@34102.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@34102.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@34102.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@34102.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@34102.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@34102.4]
  input          io_memStreams_stores_0_data_ready, // @[:@34102.4]
  output         io_memStreams_stores_0_data_valid, // @[:@34102.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@34102.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@34102.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@34102.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@34102.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@34102.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@34102.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@34102.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@34102.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@34102.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@34102.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@34102.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@34102.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@34102.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@34102.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@34102.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@34102.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@34102.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@34102.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@34102.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@34102.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@34102.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@34102.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@34102.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@34102.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@34102.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@34102.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@34102.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@34102.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@34102.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@34102.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@34102.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@34102.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@34102.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@34102.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@34102.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@34102.4]
  output         io_heap_0_req_valid, // @[:@34102.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@34102.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@34102.4]
  input          io_heap_0_resp_valid, // @[:@34102.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@34102.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@34102.4]
  input  [63:0]  io_argIns_0, // @[:@34102.4]
  input  [63:0]  io_argIns_1, // @[:@34102.4]
  input          io_argOuts_0_port_ready, // @[:@34102.4]
  output         io_argOuts_0_port_valid, // @[:@34102.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@34102.4]
  input  [63:0]  io_argOuts_0_echo // @[:@34102.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@34250.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@34250.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@34250.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@34250.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34268.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34268.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34268.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34268.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34268.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@34277.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@34277.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@34277.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@34277.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@34277.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@34277.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@34316.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34348.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34348.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34348.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34348.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34348.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x444_ready; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x444_valid; // @[sm_RootController.scala 91:24:@34410.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x444_bits_addr; // @[sm_RootController.scala 91:24:@34410.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x444_bits_size; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x445_ready; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x445_valid; // @[sm_RootController.scala 91:24:@34410.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x445_bits_wdata_0; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x445_bits_wstrb; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x241_TVALID; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x241_TREADY; // @[sm_RootController.scala 91:24:@34410.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x241_TDATA; // @[sm_RootController.scala 91:24:@34410.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x241_TID; // @[sm_RootController.scala 91:24:@34410.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x241_TDEST; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x446_ready; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x446_valid; // @[sm_RootController.scala 91:24:@34410.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x239_outdram_number; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x242_TVALID; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_in_x242_TREADY; // @[sm_RootController.scala 91:24:@34410.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x242_TDATA; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@34410.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@34410.4]
  wire  _T_599; // @[package.scala 96:25:@34273.4 package.scala 96:25:@34274.4]
  wire  _T_664; // @[Main.scala 46:50:@34344.4]
  wire  _T_665; // @[Main.scala 46:59:@34345.4]
  wire  _T_677; // @[package.scala 100:49:@34365.4]
  reg  _T_680; // @[package.scala 48:56:@34366.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@34250.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34268.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@34277.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@34316.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34348.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@34410.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x444_ready(RootController_kernelRootController_concrete1_io_in_x444_ready),
    .io_in_x444_valid(RootController_kernelRootController_concrete1_io_in_x444_valid),
    .io_in_x444_bits_addr(RootController_kernelRootController_concrete1_io_in_x444_bits_addr),
    .io_in_x444_bits_size(RootController_kernelRootController_concrete1_io_in_x444_bits_size),
    .io_in_x445_ready(RootController_kernelRootController_concrete1_io_in_x445_ready),
    .io_in_x445_valid(RootController_kernelRootController_concrete1_io_in_x445_valid),
    .io_in_x445_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x445_bits_wdata_0),
    .io_in_x445_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x445_bits_wstrb),
    .io_in_x241_TVALID(RootController_kernelRootController_concrete1_io_in_x241_TVALID),
    .io_in_x241_TREADY(RootController_kernelRootController_concrete1_io_in_x241_TREADY),
    .io_in_x241_TDATA(RootController_kernelRootController_concrete1_io_in_x241_TDATA),
    .io_in_x241_TID(RootController_kernelRootController_concrete1_io_in_x241_TID),
    .io_in_x241_TDEST(RootController_kernelRootController_concrete1_io_in_x241_TDEST),
    .io_in_x446_ready(RootController_kernelRootController_concrete1_io_in_x446_ready),
    .io_in_x446_valid(RootController_kernelRootController_concrete1_io_in_x446_valid),
    .io_in_x239_outdram_number(RootController_kernelRootController_concrete1_io_in_x239_outdram_number),
    .io_in_x242_TVALID(RootController_kernelRootController_concrete1_io_in_x242_TVALID),
    .io_in_x242_TREADY(RootController_kernelRootController_concrete1_io_in_x242_TREADY),
    .io_in_x242_TDATA(RootController_kernelRootController_concrete1_io_in_x242_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@34273.4 package.scala 96:25:@34274.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@34344.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@34345.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@34365.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@34364.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x444_valid; // @[sm_RootController.scala 60:23:@34473.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x444_bits_addr; // @[sm_RootController.scala 60:23:@34472.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x444_bits_size; // @[sm_RootController.scala 60:23:@34471.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x445_valid; // @[sm_RootController.scala 61:23:@34477.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x445_bits_wdata_0; // @[sm_RootController.scala 61:23:@34476.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x445_bits_wstrb; // @[sm_RootController.scala 61:23:@34475.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x446_ready; // @[sm_RootController.scala 63:23:@34490.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x241_TREADY; // @[sm_RootController.scala 62:23:@34486.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x242_TVALID; // @[sm_RootController.scala 65:23:@34500.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x242_TDATA; // @[sm_RootController.scala 65:23:@34498.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 65:23:@34497.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 65:23:@34496.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 65:23:@34495.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 65:23:@34494.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 65:23:@34493.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 65:23:@34492.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@34251.4]
  assign SingleCounter_reset = reset; // @[:@34252.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@34266.4]
  assign RetimeWrapper_clock = clock; // @[:@34269.4]
  assign RetimeWrapper_reset = reset; // @[:@34270.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34272.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@34271.4]
  assign SRFF_clock = clock; // @[:@34278.4]
  assign SRFF_reset = reset; // @[:@34279.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@34528.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@34362.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@34363.4]
  assign RootController_sm_clock = clock; // @[:@34317.4]
  assign RootController_sm_reset = reset; // @[:@34318.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@34361.4 SpatialBlocks.scala 140:18:@34395.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@34389.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@34369.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@34357.4 SpatialBlocks.scala 142:21:@34397.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@34386.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34349.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34350.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34352.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@34351.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@34411.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@34412.4]
  assign RootController_kernelRootController_concrete1_io_in_x444_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 60:23:@34474.4]
  assign RootController_kernelRootController_concrete1_io_in_x445_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 61:23:@34478.4]
  assign RootController_kernelRootController_concrete1_io_in_x241_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 62:23:@34487.4]
  assign RootController_kernelRootController_concrete1_io_in_x241_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 62:23:@34485.4]
  assign RootController_kernelRootController_concrete1_io_in_x241_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 62:23:@34481.4]
  assign RootController_kernelRootController_concrete1_io_in_x241_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 62:23:@34480.4]
  assign RootController_kernelRootController_concrete1_io_in_x446_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 63:23:@34489.4]
  assign RootController_kernelRootController_concrete1_io_in_x239_outdram_number = io_argIns_1; // @[sm_RootController.scala 64:31:@34491.4]
  assign RootController_kernelRootController_concrete1_io_in_x242_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 65:23:@34499.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@34509.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@34507.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@34501.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@34530.2]
  input        clock, // @[:@34531.4]
  input        reset, // @[:@34532.4]
  input        io_enable, // @[:@34533.4]
  output [5:0] io_out, // @[:@34533.4]
  output [5:0] io_next // @[:@34533.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@34535.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@34536.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@34537.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@34542.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@34536.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@34537.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@34542.6]
  assign io_out = count; // @[Counter.scala 25:10:@34545.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@34546.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_17( // @[:@34582.2]
  input         clock, // @[:@34583.4]
  input         reset, // @[:@34584.4]
  input  [5:0]  io_raddr, // @[:@34585.4]
  input         io_wen, // @[:@34585.4]
  input  [5:0]  io_waddr, // @[:@34585.4]
  input  [63:0] io_wdata_addr, // @[:@34585.4]
  input  [31:0] io_wdata_size, // @[:@34585.4]
  output [63:0] io_rdata_addr, // @[:@34585.4]
  output [31:0] io_rdata_size // @[:@34585.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@34587.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@34587.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@34587.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@34587.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@34587.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@34587.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@34587.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@34587.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@34587.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@34601.4]
  wire  _T_20; // @[SRAM.scala 182:49:@34606.4]
  wire  _T_21; // @[SRAM.scala 182:37:@34607.4]
  reg  _T_24; // @[SRAM.scala 182:29:@34608.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@34611.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@34613.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@34587.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@34601.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@34606.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@34607.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@34613.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@34622.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@34621.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@34602.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@34603.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@34599.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@34605.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@34604.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@34600.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@34598.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@34597.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@34624.2]
  input         clock, // @[:@34625.4]
  input         reset, // @[:@34626.4]
  output        io_in_ready, // @[:@34627.4]
  input         io_in_valid, // @[:@34627.4]
  input  [63:0] io_in_bits_addr, // @[:@34627.4]
  input  [31:0] io_in_bits_size, // @[:@34627.4]
  input         io_out_ready, // @[:@34627.4]
  output        io_out_valid, // @[:@34627.4]
  output [63:0] io_out_bits_addr, // @[:@34627.4]
  output [31:0] io_out_bits_size // @[:@34627.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@35023.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@35023.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@35023.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@35023.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@35023.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@35033.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@35033.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@35033.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@35033.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@35033.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@35048.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@35048.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@35048.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@35048.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@35048.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@35048.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@35048.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@35048.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@35048.4]
  wire  writeEn; // @[FIFO.scala 30:29:@35021.4]
  wire  readEn; // @[FIFO.scala 31:29:@35022.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@35043.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@35044.4]
  wire  _T_824; // @[FIFO.scala 45:27:@35045.4]
  wire  empty; // @[FIFO.scala 45:24:@35046.4]
  wire  full; // @[FIFO.scala 46:23:@35047.4]
  wire  _T_827; // @[FIFO.scala 83:17:@35060.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@35061.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@35023.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@35033.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_17 SRAM ( // @[FIFO.scala 73:19:@35048.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@35021.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@35022.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@35044.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@35045.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@35046.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@35047.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@35060.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@35061.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@35067.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@35065.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@35058.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@35057.4]
  assign enqCounter_clock = clock; // @[:@35024.4]
  assign enqCounter_reset = reset; // @[:@35025.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@35031.4]
  assign deqCounter_clock = clock; // @[:@35034.4]
  assign deqCounter_reset = reset; // @[:@35035.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@35041.4]
  assign SRAM_clock = clock; // @[:@35049.4]
  assign SRAM_reset = reset; // @[:@35050.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@35052.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@35053.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@35054.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@35056.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@35055.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@35069.2]
  input        clock, // @[:@35070.4]
  input        reset, // @[:@35071.4]
  input        io_enable, // @[:@35072.4]
  output [3:0] io_out // @[:@35072.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@35074.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@35075.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@35076.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@35081.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@35075.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@35076.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@35081.6]
  assign io_out = count; // @[Counter.scala 25:10:@35084.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@35105.2]
  input        clock, // @[:@35106.4]
  input        reset, // @[:@35107.4]
  input        io_reset, // @[:@35108.4]
  input        io_enable, // @[:@35108.4]
  input  [1:0] io_stride, // @[:@35108.4]
  output [1:0] io_out, // @[:@35108.4]
  output [1:0] io_next // @[:@35108.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@35110.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@35111.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@35112.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@35117.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@35113.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@35111.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@35112.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@35117.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@35113.4]
  assign io_out = count; // @[Counter.scala 25:10:@35120.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@35121.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_18( // @[:@35157.2]
  input         clock, // @[:@35158.4]
  input         reset, // @[:@35159.4]
  input  [1:0]  io_raddr, // @[:@35160.4]
  input         io_wen, // @[:@35160.4]
  input  [1:0]  io_waddr, // @[:@35160.4]
  input  [31:0] io_wdata, // @[:@35160.4]
  output [31:0] io_rdata, // @[:@35160.4]
  input         io_backpressure // @[:@35160.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@35162.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@35162.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@35162.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@35162.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@35162.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@35162.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@35162.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@35162.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@35162.4]
  wire  _T_19; // @[SRAM.scala 182:49:@35180.4]
  wire  _T_20; // @[SRAM.scala 182:37:@35181.4]
  reg  _T_23; // @[SRAM.scala 182:29:@35182.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@35184.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@35162.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@35180.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@35181.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@35189.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@35176.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@35177.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@35174.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@35179.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@35178.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@35175.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@35173.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@35172.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@35191.2]
  input         clock, // @[:@35192.4]
  input         reset, // @[:@35193.4]
  output        io_in_ready, // @[:@35194.4]
  input         io_in_valid, // @[:@35194.4]
  input  [31:0] io_in_bits, // @[:@35194.4]
  input         io_out_ready, // @[:@35194.4]
  output        io_out_valid, // @[:@35194.4]
  output [31:0] io_out_bits // @[:@35194.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@35220.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@35220.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@35220.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@35220.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@35220.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@35220.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@35220.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@35230.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@35230.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@35230.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@35230.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@35230.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@35230.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@35230.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@35245.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@35245.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@35245.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@35245.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@35245.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@35245.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@35245.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@35245.4]
  wire  writeEn; // @[FIFO.scala 30:29:@35218.4]
  wire  readEn; // @[FIFO.scala 31:29:@35219.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@35240.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@35241.4]
  wire  _T_104; // @[FIFO.scala 45:27:@35242.4]
  wire  empty; // @[FIFO.scala 45:24:@35243.4]
  wire  full; // @[FIFO.scala 46:23:@35244.4]
  wire  _T_107; // @[FIFO.scala 83:17:@35255.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@35256.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@35220.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@35230.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_18 SRAM ( // @[FIFO.scala 73:19:@35245.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@35218.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@35219.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@35241.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@35242.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@35243.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@35244.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@35255.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@35256.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@35262.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@35260.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@35253.4]
  assign enqCounter_clock = clock; // @[:@35221.4]
  assign enqCounter_reset = reset; // @[:@35222.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@35228.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@35229.4]
  assign deqCounter_clock = clock; // @[:@35231.4]
  assign deqCounter_reset = reset; // @[:@35232.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@35238.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@35239.4]
  assign SRAM_clock = clock; // @[:@35246.4]
  assign SRAM_reset = reset; // @[:@35247.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@35249.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@35250.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@35251.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@35252.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@35254.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@37649.2]
  input         clock, // @[:@37650.4]
  input         reset, // @[:@37651.4]
  output        io_in_ready, // @[:@37652.4]
  input         io_in_valid, // @[:@37652.4]
  input  [31:0] io_in_bits_0, // @[:@37652.4]
  input         io_out_ready, // @[:@37652.4]
  output        io_out_valid, // @[:@37652.4]
  output [31:0] io_out_bits_0, // @[:@37652.4]
  output [31:0] io_out_bits_1, // @[:@37652.4]
  output [31:0] io_out_bits_2, // @[:@37652.4]
  output [31:0] io_out_bits_3, // @[:@37652.4]
  output [31:0] io_out_bits_4, // @[:@37652.4]
  output [31:0] io_out_bits_5, // @[:@37652.4]
  output [31:0] io_out_bits_6, // @[:@37652.4]
  output [31:0] io_out_bits_7, // @[:@37652.4]
  output [31:0] io_out_bits_8, // @[:@37652.4]
  output [31:0] io_out_bits_9, // @[:@37652.4]
  output [31:0] io_out_bits_10, // @[:@37652.4]
  output [31:0] io_out_bits_11, // @[:@37652.4]
  output [31:0] io_out_bits_12, // @[:@37652.4]
  output [31:0] io_out_bits_13, // @[:@37652.4]
  output [31:0] io_out_bits_14, // @[:@37652.4]
  output [31:0] io_out_bits_15 // @[:@37652.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@37656.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@37656.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@37656.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@37656.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@37667.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@37667.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@37667.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@37667.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@37680.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@37680.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@37680.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@37680.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@37680.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@37680.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@37680.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@37680.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@37715.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@37715.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@37715.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@37715.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@37715.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@37715.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@37715.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@37715.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@37750.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@37750.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@37750.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@37750.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@37750.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@37750.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@37750.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@37750.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@37785.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@37785.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@37785.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@37785.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@37785.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@37785.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@37785.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@37785.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@37820.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@37820.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@37820.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@37820.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@37820.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@37820.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@37820.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@37820.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@37855.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@37855.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@37855.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@37855.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@37855.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@37855.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@37855.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@37855.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@37890.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@37890.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@37890.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@37890.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@37890.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@37890.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@37890.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@37890.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@37925.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@37925.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@37925.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@37925.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@37925.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@37925.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@37925.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@37925.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@37960.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@37960.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@37960.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@37960.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@37960.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@37960.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@37960.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@37960.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@37995.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@37995.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@37995.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@37995.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@37995.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@37995.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@37995.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@37995.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@38030.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@38030.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@38030.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@38030.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@38030.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@38030.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@38030.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@38030.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@38065.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@38065.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@38065.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@38065.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@38065.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@38065.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@38065.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@38065.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@38100.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@38100.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@38100.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@38100.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@38100.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@38100.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@38100.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@38100.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@38135.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@38135.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@38135.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@38135.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@38135.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@38135.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@38135.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@38135.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@38170.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@38170.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@38170.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@38170.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@38170.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@38170.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@38170.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@38170.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@38205.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@38205.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@38205.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@38205.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@38205.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@38205.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@38205.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@38205.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@37655.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@37678.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@37705.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@37740.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@37775.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@37810.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@37845.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@37880.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@37915.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@37950.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@37985.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@38020.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@38055.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@38090.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@38125.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@38160.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@38195.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@38230.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38241.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38242.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38243.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38244.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38245.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38246.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38247.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38248.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38249.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38250.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38251.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38252.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38253.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38254.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38255.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@38272.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38256.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@38291.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@38292.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@38293.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@38294.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@38295.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@38296.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@38297.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@38298.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@38299.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@38300.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@38301.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@38302.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@38303.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@38304.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@37656.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@37667.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@37680.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@37715.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@37750.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@37785.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@37820.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@37855.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@37890.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@37925.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@37960.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@37995.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@38030.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@38065.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@38100.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@38135.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@38170.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@38205.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@37655.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@37678.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@37705.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@37740.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@37775.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@37810.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@37845.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@37880.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@37915.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@37950.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@37985.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@38020.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@38055.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@38090.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@38125.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@38160.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@38195.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@38230.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38241.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38242.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38243.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38244.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38245.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38246.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38247.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38248.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38249.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38250.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38251.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38252.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38253.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38254.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38255.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@38272.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@38240.4 FIFOVec.scala 49:42:@38256.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@38291.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@38292.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@38293.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@38294.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@38295.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@38296.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@38297.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@38298.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@38299.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@38300.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@38301.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@38302.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@38303.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@38304.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@38273.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@38307.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@38615.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@38616.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@38617.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@38618.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@38619.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@38620.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@38621.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@38622.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@38623.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@38624.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@38625.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@38626.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@38627.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@38628.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@38629.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@38630.4]
  assign enqCounter_clock = clock; // @[:@37657.4]
  assign enqCounter_reset = reset; // @[:@37658.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@37665.4]
  assign deqCounter_clock = clock; // @[:@37668.4]
  assign deqCounter_reset = reset; // @[:@37669.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@37676.4]
  assign fifos_0_clock = clock; // @[:@37681.4]
  assign fifos_0_reset = reset; // @[:@37682.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@37708.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37710.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37714.4]
  assign fifos_1_clock = clock; // @[:@37716.4]
  assign fifos_1_reset = reset; // @[:@37717.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@37743.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37745.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37749.4]
  assign fifos_2_clock = clock; // @[:@37751.4]
  assign fifos_2_reset = reset; // @[:@37752.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@37778.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37780.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37784.4]
  assign fifos_3_clock = clock; // @[:@37786.4]
  assign fifos_3_reset = reset; // @[:@37787.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@37813.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37815.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37819.4]
  assign fifos_4_clock = clock; // @[:@37821.4]
  assign fifos_4_reset = reset; // @[:@37822.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@37848.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37850.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37854.4]
  assign fifos_5_clock = clock; // @[:@37856.4]
  assign fifos_5_reset = reset; // @[:@37857.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@37883.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37885.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37889.4]
  assign fifos_6_clock = clock; // @[:@37891.4]
  assign fifos_6_reset = reset; // @[:@37892.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@37918.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37920.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37924.4]
  assign fifos_7_clock = clock; // @[:@37926.4]
  assign fifos_7_reset = reset; // @[:@37927.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@37953.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37955.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37959.4]
  assign fifos_8_clock = clock; // @[:@37961.4]
  assign fifos_8_reset = reset; // @[:@37962.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@37988.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37990.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37994.4]
  assign fifos_9_clock = clock; // @[:@37996.4]
  assign fifos_9_reset = reset; // @[:@37997.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@38023.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38025.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38029.4]
  assign fifos_10_clock = clock; // @[:@38031.4]
  assign fifos_10_reset = reset; // @[:@38032.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@38058.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38060.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38064.4]
  assign fifos_11_clock = clock; // @[:@38066.4]
  assign fifos_11_reset = reset; // @[:@38067.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@38093.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38095.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38099.4]
  assign fifos_12_clock = clock; // @[:@38101.4]
  assign fifos_12_reset = reset; // @[:@38102.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@38128.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38130.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38134.4]
  assign fifos_13_clock = clock; // @[:@38136.4]
  assign fifos_13_reset = reset; // @[:@38137.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@38163.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38165.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38169.4]
  assign fifos_14_clock = clock; // @[:@38171.4]
  assign fifos_14_reset = reset; // @[:@38172.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@38198.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38200.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38204.4]
  assign fifos_15_clock = clock; // @[:@38206.4]
  assign fifos_15_reset = reset; // @[:@38207.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@38233.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38235.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38239.4]
endmodule
module FFRAM( // @[:@38704.2]
  input        clock, // @[:@38705.4]
  input        reset, // @[:@38706.4]
  input  [1:0] io_raddr, // @[:@38707.4]
  input        io_wen, // @[:@38707.4]
  input  [1:0] io_waddr, // @[:@38707.4]
  input        io_wdata, // @[:@38707.4]
  output       io_rdata, // @[:@38707.4]
  input        io_banks_0_wdata_valid, // @[:@38707.4]
  input        io_banks_0_wdata_bits, // @[:@38707.4]
  input        io_banks_1_wdata_valid, // @[:@38707.4]
  input        io_banks_1_wdata_bits, // @[:@38707.4]
  input        io_banks_2_wdata_valid, // @[:@38707.4]
  input        io_banks_2_wdata_bits, // @[:@38707.4]
  input        io_banks_3_wdata_valid, // @[:@38707.4]
  input        io_banks_3_wdata_bits // @[:@38707.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@38711.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@38712.4]
  wire  _T_89; // @[SRAM.scala 148:25:@38713.4]
  wire  _T_90; // @[SRAM.scala 148:15:@38714.4]
  wire  _T_91; // @[SRAM.scala 149:15:@38716.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@38715.4]
  reg  regs_1; // @[SRAM.scala 145:20:@38722.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@38723.4]
  wire  _T_98; // @[SRAM.scala 148:25:@38724.4]
  wire  _T_99; // @[SRAM.scala 148:15:@38725.4]
  wire  _T_100; // @[SRAM.scala 149:15:@38727.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@38726.4]
  reg  regs_2; // @[SRAM.scala 145:20:@38733.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@38734.4]
  wire  _T_107; // @[SRAM.scala 148:25:@38735.4]
  wire  _T_108; // @[SRAM.scala 148:15:@38736.4]
  wire  _T_109; // @[SRAM.scala 149:15:@38738.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@38737.4]
  reg  regs_3; // @[SRAM.scala 145:20:@38744.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@38745.4]
  wire  _T_116; // @[SRAM.scala 148:25:@38746.4]
  wire  _T_117; // @[SRAM.scala 148:15:@38747.4]
  wire  _T_118; // @[SRAM.scala 149:15:@38749.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@38748.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@38758.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@38758.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@38712.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@38713.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@38714.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38716.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@38715.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@38723.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@38724.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@38725.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38727.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@38726.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@38734.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@38735.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@38736.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38738.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@38737.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@38745.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@38746.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@38747.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38749.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@38748.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@38758.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@38758.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@38758.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@38760.2]
  input   clock, // @[:@38761.4]
  input   reset, // @[:@38762.4]
  output  io_in_ready, // @[:@38763.4]
  input   io_in_valid, // @[:@38763.4]
  input   io_in_bits, // @[:@38763.4]
  input   io_out_ready, // @[:@38763.4]
  output  io_out_valid, // @[:@38763.4]
  output  io_out_bits // @[:@38763.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@38789.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@38789.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@38789.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@38789.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@38789.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@38789.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@38789.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@38799.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@38799.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@38799.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@38799.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@38799.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@38799.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@38799.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@38814.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@38814.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@38814.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@38814.4]
  wire  writeEn; // @[FIFO.scala 30:29:@38787.4]
  wire  readEn; // @[FIFO.scala 31:29:@38788.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@38809.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@38810.4]
  wire  _T_104; // @[FIFO.scala 45:27:@38811.4]
  wire  empty; // @[FIFO.scala 45:24:@38812.4]
  wire  full; // @[FIFO.scala 46:23:@38813.4]
  wire  _T_157; // @[FIFO.scala 83:17:@38900.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@38901.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@38789.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@38799.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@38814.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@38787.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@38788.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@38810.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@38811.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@38812.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@38813.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@38900.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@38901.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@38907.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@38905.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@38839.4]
  assign enqCounter_clock = clock; // @[:@38790.4]
  assign enqCounter_reset = reset; // @[:@38791.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@38797.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@38798.4]
  assign deqCounter_clock = clock; // @[:@38800.4]
  assign deqCounter_reset = reset; // @[:@38801.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@38807.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@38808.4]
  assign FFRAM_clock = clock; // @[:@38815.4]
  assign FFRAM_reset = reset; // @[:@38816.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@38835.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@38836.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@38837.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@38838.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38841.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38840.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38844.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38843.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38847.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38846.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38850.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38849.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@42524.2]
  input   clock, // @[:@42525.4]
  input   reset, // @[:@42526.4]
  output  io_in_ready, // @[:@42527.4]
  input   io_in_valid, // @[:@42527.4]
  input   io_in_bits_0, // @[:@42527.4]
  input   io_out_ready, // @[:@42527.4]
  output  io_out_valid, // @[:@42527.4]
  output  io_out_bits_0, // @[:@42527.4]
  output  io_out_bits_1, // @[:@42527.4]
  output  io_out_bits_2, // @[:@42527.4]
  output  io_out_bits_3, // @[:@42527.4]
  output  io_out_bits_4, // @[:@42527.4]
  output  io_out_bits_5, // @[:@42527.4]
  output  io_out_bits_6, // @[:@42527.4]
  output  io_out_bits_7, // @[:@42527.4]
  output  io_out_bits_8, // @[:@42527.4]
  output  io_out_bits_9, // @[:@42527.4]
  output  io_out_bits_10, // @[:@42527.4]
  output  io_out_bits_11, // @[:@42527.4]
  output  io_out_bits_12, // @[:@42527.4]
  output  io_out_bits_13, // @[:@42527.4]
  output  io_out_bits_14, // @[:@42527.4]
  output  io_out_bits_15 // @[:@42527.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@42531.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@42531.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@42531.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@42531.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@42542.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@42542.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@42542.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@42542.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@42555.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@42590.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@42625.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@42660.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@42695.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@42730.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@42765.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@42800.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@42835.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@42870.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@42905.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@42940.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@42975.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@43010.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@43045.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@43080.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@43080.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@43080.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@43080.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@43080.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@43080.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@43080.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@43080.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@42530.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@42553.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@42580.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@42615.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@42650.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@42685.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@42720.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@42755.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@42790.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@42825.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@42860.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@42895.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@42930.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@42965.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@43000.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@43035.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@43070.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@43105.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43116.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43117.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43118.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43119.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43120.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43121.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43122.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43123.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43124.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43125.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43126.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43127.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43128.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43129.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43130.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@43147.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43131.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@43166.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@43167.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@43168.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@43169.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@43170.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@43171.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@43172.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@43173.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@43174.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@43175.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@43176.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@43177.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@43178.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@43179.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@42531.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@42542.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@42555.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@42590.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@42625.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@42660.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@42695.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@42730.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@42765.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@42800.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@42835.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@42870.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@42905.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@42940.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@42975.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@43010.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@43045.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@43080.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@42530.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@42553.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@42580.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@42615.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@42650.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@42685.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@42720.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@42755.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@42790.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@42825.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@42860.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@42895.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@42930.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@42965.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@43000.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@43035.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@43070.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@43105.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43116.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43117.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43118.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43119.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43120.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43121.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43122.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43123.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43124.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43125.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43126.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43127.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43128.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43129.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43130.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@43147.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@43115.4 FIFOVec.scala 49:42:@43131.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@43166.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@43167.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@43168.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@43169.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@43170.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@43171.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@43172.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@43173.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@43174.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@43175.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@43176.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@43177.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@43178.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@43179.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@43148.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@43182.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@43490.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@43491.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@43492.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@43493.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@43494.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@43495.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@43496.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@43497.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@43498.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@43499.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@43500.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@43501.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@43502.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@43503.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@43504.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@43505.4]
  assign enqCounter_clock = clock; // @[:@42532.4]
  assign enqCounter_reset = reset; // @[:@42533.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@42540.4]
  assign deqCounter_clock = clock; // @[:@42543.4]
  assign deqCounter_reset = reset; // @[:@42544.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@42551.4]
  assign fifos_0_clock = clock; // @[:@42556.4]
  assign fifos_0_reset = reset; // @[:@42557.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@42583.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42585.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42589.4]
  assign fifos_1_clock = clock; // @[:@42591.4]
  assign fifos_1_reset = reset; // @[:@42592.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@42618.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42620.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42624.4]
  assign fifos_2_clock = clock; // @[:@42626.4]
  assign fifos_2_reset = reset; // @[:@42627.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@42653.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42655.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42659.4]
  assign fifos_3_clock = clock; // @[:@42661.4]
  assign fifos_3_reset = reset; // @[:@42662.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@42688.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42690.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42694.4]
  assign fifos_4_clock = clock; // @[:@42696.4]
  assign fifos_4_reset = reset; // @[:@42697.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@42723.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42725.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42729.4]
  assign fifos_5_clock = clock; // @[:@42731.4]
  assign fifos_5_reset = reset; // @[:@42732.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@42758.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42760.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42764.4]
  assign fifos_6_clock = clock; // @[:@42766.4]
  assign fifos_6_reset = reset; // @[:@42767.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@42793.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42795.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42799.4]
  assign fifos_7_clock = clock; // @[:@42801.4]
  assign fifos_7_reset = reset; // @[:@42802.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@42828.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42830.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42834.4]
  assign fifos_8_clock = clock; // @[:@42836.4]
  assign fifos_8_reset = reset; // @[:@42837.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@42863.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42865.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42869.4]
  assign fifos_9_clock = clock; // @[:@42871.4]
  assign fifos_9_reset = reset; // @[:@42872.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@42898.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42900.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42904.4]
  assign fifos_10_clock = clock; // @[:@42906.4]
  assign fifos_10_reset = reset; // @[:@42907.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@42933.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42935.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42939.4]
  assign fifos_11_clock = clock; // @[:@42941.4]
  assign fifos_11_reset = reset; // @[:@42942.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@42968.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42970.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42974.4]
  assign fifos_12_clock = clock; // @[:@42976.4]
  assign fifos_12_reset = reset; // @[:@42977.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@43003.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43005.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43009.4]
  assign fifos_13_clock = clock; // @[:@43011.4]
  assign fifos_13_reset = reset; // @[:@43012.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@43038.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43040.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43044.4]
  assign fifos_14_clock = clock; // @[:@43046.4]
  assign fifos_14_reset = reset; // @[:@43047.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@43073.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43075.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43079.4]
  assign fifos_15_clock = clock; // @[:@43081.4]
  assign fifos_15_reset = reset; // @[:@43082.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@43108.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43110.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43114.4]
endmodule
module FIFOWidthConvert( // @[:@43507.2]
  input         clock, // @[:@43508.4]
  input         reset, // @[:@43509.4]
  output        io_in_ready, // @[:@43510.4]
  input         io_in_valid, // @[:@43510.4]
  input  [31:0] io_in_bits_data_0, // @[:@43510.4]
  input         io_in_bits_strobe, // @[:@43510.4]
  input         io_out_ready, // @[:@43510.4]
  output        io_out_valid, // @[:@43510.4]
  output [31:0] io_out_bits_data_0, // @[:@43510.4]
  output [31:0] io_out_bits_data_1, // @[:@43510.4]
  output [31:0] io_out_bits_data_2, // @[:@43510.4]
  output [31:0] io_out_bits_data_3, // @[:@43510.4]
  output [31:0] io_out_bits_data_4, // @[:@43510.4]
  output [31:0] io_out_bits_data_5, // @[:@43510.4]
  output [31:0] io_out_bits_data_6, // @[:@43510.4]
  output [31:0] io_out_bits_data_7, // @[:@43510.4]
  output [31:0] io_out_bits_data_8, // @[:@43510.4]
  output [31:0] io_out_bits_data_9, // @[:@43510.4]
  output [31:0] io_out_bits_data_10, // @[:@43510.4]
  output [31:0] io_out_bits_data_11, // @[:@43510.4]
  output [31:0] io_out_bits_data_12, // @[:@43510.4]
  output [31:0] io_out_bits_data_13, // @[:@43510.4]
  output [31:0] io_out_bits_data_14, // @[:@43510.4]
  output [31:0] io_out_bits_data_15, // @[:@43510.4]
  output [63:0] io_out_bits_strobe // @[:@43510.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@43512.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@43553.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@43612.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@43618.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@43676.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@43682.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@43683.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@43687.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@43691.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@43695.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@43699.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@43703.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@43707.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@43711.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@43715.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@43719.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@43723.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@43727.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@43731.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@43735.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@43739.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@43743.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@43820.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@43829.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@43838.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@43847.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@43856.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@43865.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@43873.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@43512.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@43553.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@43612.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@43618.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@43676.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@43682.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@43683.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@43687.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@43691.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@43695.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@43699.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@43703.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@43707.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@43711.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@43715.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@43719.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@43723.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@43727.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@43731.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@43735.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@43739.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@43743.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@43820.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@43829.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@43838.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@43847.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@43856.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@43865.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@43873.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@43602.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@43603.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@43652.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@43653.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@43654.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@43655.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@43656.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@43657.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@43658.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@43659.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@43660.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@43661.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@43662.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@43663.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@43664.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@43665.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@43666.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@43667.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@43875.4]
  assign FIFOVec_clock = clock; // @[:@43513.4]
  assign FIFOVec_reset = reset; // @[:@43514.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@43599.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@43598.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@43876.4]
  assign FIFOVec_1_clock = clock; // @[:@43554.4]
  assign FIFOVec_1_reset = reset; // @[:@43555.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@43601.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@43600.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@43877.4]
endmodule
module FFRAM_16( // @[:@43915.2]
  input        clock, // @[:@43916.4]
  input        reset, // @[:@43917.4]
  input  [5:0] io_raddr, // @[:@43918.4]
  input        io_wen, // @[:@43918.4]
  input  [5:0] io_waddr, // @[:@43918.4]
  input        io_wdata, // @[:@43918.4]
  output       io_rdata, // @[:@43918.4]
  input        io_banks_0_wdata_valid, // @[:@43918.4]
  input        io_banks_0_wdata_bits, // @[:@43918.4]
  input        io_banks_1_wdata_valid, // @[:@43918.4]
  input        io_banks_1_wdata_bits, // @[:@43918.4]
  input        io_banks_2_wdata_valid, // @[:@43918.4]
  input        io_banks_2_wdata_bits, // @[:@43918.4]
  input        io_banks_3_wdata_valid, // @[:@43918.4]
  input        io_banks_3_wdata_bits, // @[:@43918.4]
  input        io_banks_4_wdata_valid, // @[:@43918.4]
  input        io_banks_4_wdata_bits, // @[:@43918.4]
  input        io_banks_5_wdata_valid, // @[:@43918.4]
  input        io_banks_5_wdata_bits, // @[:@43918.4]
  input        io_banks_6_wdata_valid, // @[:@43918.4]
  input        io_banks_6_wdata_bits, // @[:@43918.4]
  input        io_banks_7_wdata_valid, // @[:@43918.4]
  input        io_banks_7_wdata_bits, // @[:@43918.4]
  input        io_banks_8_wdata_valid, // @[:@43918.4]
  input        io_banks_8_wdata_bits, // @[:@43918.4]
  input        io_banks_9_wdata_valid, // @[:@43918.4]
  input        io_banks_9_wdata_bits, // @[:@43918.4]
  input        io_banks_10_wdata_valid, // @[:@43918.4]
  input        io_banks_10_wdata_bits, // @[:@43918.4]
  input        io_banks_11_wdata_valid, // @[:@43918.4]
  input        io_banks_11_wdata_bits, // @[:@43918.4]
  input        io_banks_12_wdata_valid, // @[:@43918.4]
  input        io_banks_12_wdata_bits, // @[:@43918.4]
  input        io_banks_13_wdata_valid, // @[:@43918.4]
  input        io_banks_13_wdata_bits, // @[:@43918.4]
  input        io_banks_14_wdata_valid, // @[:@43918.4]
  input        io_banks_14_wdata_bits, // @[:@43918.4]
  input        io_banks_15_wdata_valid, // @[:@43918.4]
  input        io_banks_15_wdata_bits, // @[:@43918.4]
  input        io_banks_16_wdata_valid, // @[:@43918.4]
  input        io_banks_16_wdata_bits, // @[:@43918.4]
  input        io_banks_17_wdata_valid, // @[:@43918.4]
  input        io_banks_17_wdata_bits, // @[:@43918.4]
  input        io_banks_18_wdata_valid, // @[:@43918.4]
  input        io_banks_18_wdata_bits, // @[:@43918.4]
  input        io_banks_19_wdata_valid, // @[:@43918.4]
  input        io_banks_19_wdata_bits, // @[:@43918.4]
  input        io_banks_20_wdata_valid, // @[:@43918.4]
  input        io_banks_20_wdata_bits, // @[:@43918.4]
  input        io_banks_21_wdata_valid, // @[:@43918.4]
  input        io_banks_21_wdata_bits, // @[:@43918.4]
  input        io_banks_22_wdata_valid, // @[:@43918.4]
  input        io_banks_22_wdata_bits, // @[:@43918.4]
  input        io_banks_23_wdata_valid, // @[:@43918.4]
  input        io_banks_23_wdata_bits, // @[:@43918.4]
  input        io_banks_24_wdata_valid, // @[:@43918.4]
  input        io_banks_24_wdata_bits, // @[:@43918.4]
  input        io_banks_25_wdata_valid, // @[:@43918.4]
  input        io_banks_25_wdata_bits, // @[:@43918.4]
  input        io_banks_26_wdata_valid, // @[:@43918.4]
  input        io_banks_26_wdata_bits, // @[:@43918.4]
  input        io_banks_27_wdata_valid, // @[:@43918.4]
  input        io_banks_27_wdata_bits, // @[:@43918.4]
  input        io_banks_28_wdata_valid, // @[:@43918.4]
  input        io_banks_28_wdata_bits, // @[:@43918.4]
  input        io_banks_29_wdata_valid, // @[:@43918.4]
  input        io_banks_29_wdata_bits, // @[:@43918.4]
  input        io_banks_30_wdata_valid, // @[:@43918.4]
  input        io_banks_30_wdata_bits, // @[:@43918.4]
  input        io_banks_31_wdata_valid, // @[:@43918.4]
  input        io_banks_31_wdata_bits, // @[:@43918.4]
  input        io_banks_32_wdata_valid, // @[:@43918.4]
  input        io_banks_32_wdata_bits, // @[:@43918.4]
  input        io_banks_33_wdata_valid, // @[:@43918.4]
  input        io_banks_33_wdata_bits, // @[:@43918.4]
  input        io_banks_34_wdata_valid, // @[:@43918.4]
  input        io_banks_34_wdata_bits, // @[:@43918.4]
  input        io_banks_35_wdata_valid, // @[:@43918.4]
  input        io_banks_35_wdata_bits, // @[:@43918.4]
  input        io_banks_36_wdata_valid, // @[:@43918.4]
  input        io_banks_36_wdata_bits, // @[:@43918.4]
  input        io_banks_37_wdata_valid, // @[:@43918.4]
  input        io_banks_37_wdata_bits, // @[:@43918.4]
  input        io_banks_38_wdata_valid, // @[:@43918.4]
  input        io_banks_38_wdata_bits, // @[:@43918.4]
  input        io_banks_39_wdata_valid, // @[:@43918.4]
  input        io_banks_39_wdata_bits, // @[:@43918.4]
  input        io_banks_40_wdata_valid, // @[:@43918.4]
  input        io_banks_40_wdata_bits, // @[:@43918.4]
  input        io_banks_41_wdata_valid, // @[:@43918.4]
  input        io_banks_41_wdata_bits, // @[:@43918.4]
  input        io_banks_42_wdata_valid, // @[:@43918.4]
  input        io_banks_42_wdata_bits, // @[:@43918.4]
  input        io_banks_43_wdata_valid, // @[:@43918.4]
  input        io_banks_43_wdata_bits, // @[:@43918.4]
  input        io_banks_44_wdata_valid, // @[:@43918.4]
  input        io_banks_44_wdata_bits, // @[:@43918.4]
  input        io_banks_45_wdata_valid, // @[:@43918.4]
  input        io_banks_45_wdata_bits, // @[:@43918.4]
  input        io_banks_46_wdata_valid, // @[:@43918.4]
  input        io_banks_46_wdata_bits, // @[:@43918.4]
  input        io_banks_47_wdata_valid, // @[:@43918.4]
  input        io_banks_47_wdata_bits, // @[:@43918.4]
  input        io_banks_48_wdata_valid, // @[:@43918.4]
  input        io_banks_48_wdata_bits, // @[:@43918.4]
  input        io_banks_49_wdata_valid, // @[:@43918.4]
  input        io_banks_49_wdata_bits, // @[:@43918.4]
  input        io_banks_50_wdata_valid, // @[:@43918.4]
  input        io_banks_50_wdata_bits, // @[:@43918.4]
  input        io_banks_51_wdata_valid, // @[:@43918.4]
  input        io_banks_51_wdata_bits, // @[:@43918.4]
  input        io_banks_52_wdata_valid, // @[:@43918.4]
  input        io_banks_52_wdata_bits, // @[:@43918.4]
  input        io_banks_53_wdata_valid, // @[:@43918.4]
  input        io_banks_53_wdata_bits, // @[:@43918.4]
  input        io_banks_54_wdata_valid, // @[:@43918.4]
  input        io_banks_54_wdata_bits, // @[:@43918.4]
  input        io_banks_55_wdata_valid, // @[:@43918.4]
  input        io_banks_55_wdata_bits, // @[:@43918.4]
  input        io_banks_56_wdata_valid, // @[:@43918.4]
  input        io_banks_56_wdata_bits, // @[:@43918.4]
  input        io_banks_57_wdata_valid, // @[:@43918.4]
  input        io_banks_57_wdata_bits, // @[:@43918.4]
  input        io_banks_58_wdata_valid, // @[:@43918.4]
  input        io_banks_58_wdata_bits, // @[:@43918.4]
  input        io_banks_59_wdata_valid, // @[:@43918.4]
  input        io_banks_59_wdata_bits, // @[:@43918.4]
  input        io_banks_60_wdata_valid, // @[:@43918.4]
  input        io_banks_60_wdata_bits, // @[:@43918.4]
  input        io_banks_61_wdata_valid, // @[:@43918.4]
  input        io_banks_61_wdata_bits, // @[:@43918.4]
  input        io_banks_62_wdata_valid, // @[:@43918.4]
  input        io_banks_62_wdata_bits, // @[:@43918.4]
  input        io_banks_63_wdata_valid, // @[:@43918.4]
  input        io_banks_63_wdata_bits // @[:@43918.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@43922.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@43923.4]
  wire  _T_689; // @[SRAM.scala 148:25:@43924.4]
  wire  _T_690; // @[SRAM.scala 148:15:@43925.4]
  wire  _T_691; // @[SRAM.scala 149:15:@43927.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@43926.4]
  reg  regs_1; // @[SRAM.scala 145:20:@43933.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@43934.4]
  wire  _T_698; // @[SRAM.scala 148:25:@43935.4]
  wire  _T_699; // @[SRAM.scala 148:15:@43936.4]
  wire  _T_700; // @[SRAM.scala 149:15:@43938.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@43937.4]
  reg  regs_2; // @[SRAM.scala 145:20:@43944.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@43945.4]
  wire  _T_707; // @[SRAM.scala 148:25:@43946.4]
  wire  _T_708; // @[SRAM.scala 148:15:@43947.4]
  wire  _T_709; // @[SRAM.scala 149:15:@43949.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@43948.4]
  reg  regs_3; // @[SRAM.scala 145:20:@43955.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@43956.4]
  wire  _T_716; // @[SRAM.scala 148:25:@43957.4]
  wire  _T_717; // @[SRAM.scala 148:15:@43958.4]
  wire  _T_718; // @[SRAM.scala 149:15:@43960.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@43959.4]
  reg  regs_4; // @[SRAM.scala 145:20:@43966.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@43967.4]
  wire  _T_725; // @[SRAM.scala 148:25:@43968.4]
  wire  _T_726; // @[SRAM.scala 148:15:@43969.4]
  wire  _T_727; // @[SRAM.scala 149:15:@43971.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@43970.4]
  reg  regs_5; // @[SRAM.scala 145:20:@43977.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@43978.4]
  wire  _T_734; // @[SRAM.scala 148:25:@43979.4]
  wire  _T_735; // @[SRAM.scala 148:15:@43980.4]
  wire  _T_736; // @[SRAM.scala 149:15:@43982.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@43981.4]
  reg  regs_6; // @[SRAM.scala 145:20:@43988.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@43989.4]
  wire  _T_743; // @[SRAM.scala 148:25:@43990.4]
  wire  _T_744; // @[SRAM.scala 148:15:@43991.4]
  wire  _T_745; // @[SRAM.scala 149:15:@43993.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@43992.4]
  reg  regs_7; // @[SRAM.scala 145:20:@43999.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@44000.4]
  wire  _T_752; // @[SRAM.scala 148:25:@44001.4]
  wire  _T_753; // @[SRAM.scala 148:15:@44002.4]
  wire  _T_754; // @[SRAM.scala 149:15:@44004.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@44003.4]
  reg  regs_8; // @[SRAM.scala 145:20:@44010.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@44011.4]
  wire  _T_761; // @[SRAM.scala 148:25:@44012.4]
  wire  _T_762; // @[SRAM.scala 148:15:@44013.4]
  wire  _T_763; // @[SRAM.scala 149:15:@44015.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@44014.4]
  reg  regs_9; // @[SRAM.scala 145:20:@44021.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@44022.4]
  wire  _T_770; // @[SRAM.scala 148:25:@44023.4]
  wire  _T_771; // @[SRAM.scala 148:15:@44024.4]
  wire  _T_772; // @[SRAM.scala 149:15:@44026.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@44025.4]
  reg  regs_10; // @[SRAM.scala 145:20:@44032.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@44033.4]
  wire  _T_779; // @[SRAM.scala 148:25:@44034.4]
  wire  _T_780; // @[SRAM.scala 148:15:@44035.4]
  wire  _T_781; // @[SRAM.scala 149:15:@44037.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@44036.4]
  reg  regs_11; // @[SRAM.scala 145:20:@44043.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@44044.4]
  wire  _T_788; // @[SRAM.scala 148:25:@44045.4]
  wire  _T_789; // @[SRAM.scala 148:15:@44046.4]
  wire  _T_790; // @[SRAM.scala 149:15:@44048.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@44047.4]
  reg  regs_12; // @[SRAM.scala 145:20:@44054.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@44055.4]
  wire  _T_797; // @[SRAM.scala 148:25:@44056.4]
  wire  _T_798; // @[SRAM.scala 148:15:@44057.4]
  wire  _T_799; // @[SRAM.scala 149:15:@44059.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@44058.4]
  reg  regs_13; // @[SRAM.scala 145:20:@44065.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@44066.4]
  wire  _T_806; // @[SRAM.scala 148:25:@44067.4]
  wire  _T_807; // @[SRAM.scala 148:15:@44068.4]
  wire  _T_808; // @[SRAM.scala 149:15:@44070.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@44069.4]
  reg  regs_14; // @[SRAM.scala 145:20:@44076.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@44077.4]
  wire  _T_815; // @[SRAM.scala 148:25:@44078.4]
  wire  _T_816; // @[SRAM.scala 148:15:@44079.4]
  wire  _T_817; // @[SRAM.scala 149:15:@44081.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@44080.4]
  reg  regs_15; // @[SRAM.scala 145:20:@44087.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@44088.4]
  wire  _T_824; // @[SRAM.scala 148:25:@44089.4]
  wire  _T_825; // @[SRAM.scala 148:15:@44090.4]
  wire  _T_826; // @[SRAM.scala 149:15:@44092.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@44091.4]
  reg  regs_16; // @[SRAM.scala 145:20:@44098.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@44099.4]
  wire  _T_833; // @[SRAM.scala 148:25:@44100.4]
  wire  _T_834; // @[SRAM.scala 148:15:@44101.4]
  wire  _T_835; // @[SRAM.scala 149:15:@44103.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@44102.4]
  reg  regs_17; // @[SRAM.scala 145:20:@44109.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@44110.4]
  wire  _T_842; // @[SRAM.scala 148:25:@44111.4]
  wire  _T_843; // @[SRAM.scala 148:15:@44112.4]
  wire  _T_844; // @[SRAM.scala 149:15:@44114.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@44113.4]
  reg  regs_18; // @[SRAM.scala 145:20:@44120.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@44121.4]
  wire  _T_851; // @[SRAM.scala 148:25:@44122.4]
  wire  _T_852; // @[SRAM.scala 148:15:@44123.4]
  wire  _T_853; // @[SRAM.scala 149:15:@44125.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@44124.4]
  reg  regs_19; // @[SRAM.scala 145:20:@44131.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@44132.4]
  wire  _T_860; // @[SRAM.scala 148:25:@44133.4]
  wire  _T_861; // @[SRAM.scala 148:15:@44134.4]
  wire  _T_862; // @[SRAM.scala 149:15:@44136.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@44135.4]
  reg  regs_20; // @[SRAM.scala 145:20:@44142.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@44143.4]
  wire  _T_869; // @[SRAM.scala 148:25:@44144.4]
  wire  _T_870; // @[SRAM.scala 148:15:@44145.4]
  wire  _T_871; // @[SRAM.scala 149:15:@44147.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@44146.4]
  reg  regs_21; // @[SRAM.scala 145:20:@44153.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@44154.4]
  wire  _T_878; // @[SRAM.scala 148:25:@44155.4]
  wire  _T_879; // @[SRAM.scala 148:15:@44156.4]
  wire  _T_880; // @[SRAM.scala 149:15:@44158.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@44157.4]
  reg  regs_22; // @[SRAM.scala 145:20:@44164.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@44165.4]
  wire  _T_887; // @[SRAM.scala 148:25:@44166.4]
  wire  _T_888; // @[SRAM.scala 148:15:@44167.4]
  wire  _T_889; // @[SRAM.scala 149:15:@44169.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@44168.4]
  reg  regs_23; // @[SRAM.scala 145:20:@44175.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@44176.4]
  wire  _T_896; // @[SRAM.scala 148:25:@44177.4]
  wire  _T_897; // @[SRAM.scala 148:15:@44178.4]
  wire  _T_898; // @[SRAM.scala 149:15:@44180.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@44179.4]
  reg  regs_24; // @[SRAM.scala 145:20:@44186.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@44187.4]
  wire  _T_905; // @[SRAM.scala 148:25:@44188.4]
  wire  _T_906; // @[SRAM.scala 148:15:@44189.4]
  wire  _T_907; // @[SRAM.scala 149:15:@44191.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@44190.4]
  reg  regs_25; // @[SRAM.scala 145:20:@44197.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@44198.4]
  wire  _T_914; // @[SRAM.scala 148:25:@44199.4]
  wire  _T_915; // @[SRAM.scala 148:15:@44200.4]
  wire  _T_916; // @[SRAM.scala 149:15:@44202.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@44201.4]
  reg  regs_26; // @[SRAM.scala 145:20:@44208.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@44209.4]
  wire  _T_923; // @[SRAM.scala 148:25:@44210.4]
  wire  _T_924; // @[SRAM.scala 148:15:@44211.4]
  wire  _T_925; // @[SRAM.scala 149:15:@44213.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@44212.4]
  reg  regs_27; // @[SRAM.scala 145:20:@44219.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@44220.4]
  wire  _T_932; // @[SRAM.scala 148:25:@44221.4]
  wire  _T_933; // @[SRAM.scala 148:15:@44222.4]
  wire  _T_934; // @[SRAM.scala 149:15:@44224.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@44223.4]
  reg  regs_28; // @[SRAM.scala 145:20:@44230.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@44231.4]
  wire  _T_941; // @[SRAM.scala 148:25:@44232.4]
  wire  _T_942; // @[SRAM.scala 148:15:@44233.4]
  wire  _T_943; // @[SRAM.scala 149:15:@44235.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@44234.4]
  reg  regs_29; // @[SRAM.scala 145:20:@44241.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@44242.4]
  wire  _T_950; // @[SRAM.scala 148:25:@44243.4]
  wire  _T_951; // @[SRAM.scala 148:15:@44244.4]
  wire  _T_952; // @[SRAM.scala 149:15:@44246.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@44245.4]
  reg  regs_30; // @[SRAM.scala 145:20:@44252.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@44253.4]
  wire  _T_959; // @[SRAM.scala 148:25:@44254.4]
  wire  _T_960; // @[SRAM.scala 148:15:@44255.4]
  wire  _T_961; // @[SRAM.scala 149:15:@44257.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@44256.4]
  reg  regs_31; // @[SRAM.scala 145:20:@44263.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@44264.4]
  wire  _T_968; // @[SRAM.scala 148:25:@44265.4]
  wire  _T_969; // @[SRAM.scala 148:15:@44266.4]
  wire  _T_970; // @[SRAM.scala 149:15:@44268.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@44267.4]
  reg  regs_32; // @[SRAM.scala 145:20:@44274.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@44275.4]
  wire  _T_977; // @[SRAM.scala 148:25:@44276.4]
  wire  _T_978; // @[SRAM.scala 148:15:@44277.4]
  wire  _T_979; // @[SRAM.scala 149:15:@44279.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@44278.4]
  reg  regs_33; // @[SRAM.scala 145:20:@44285.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@44286.4]
  wire  _T_986; // @[SRAM.scala 148:25:@44287.4]
  wire  _T_987; // @[SRAM.scala 148:15:@44288.4]
  wire  _T_988; // @[SRAM.scala 149:15:@44290.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@44289.4]
  reg  regs_34; // @[SRAM.scala 145:20:@44296.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@44297.4]
  wire  _T_995; // @[SRAM.scala 148:25:@44298.4]
  wire  _T_996; // @[SRAM.scala 148:15:@44299.4]
  wire  _T_997; // @[SRAM.scala 149:15:@44301.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@44300.4]
  reg  regs_35; // @[SRAM.scala 145:20:@44307.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@44308.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@44309.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@44310.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@44312.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@44311.4]
  reg  regs_36; // @[SRAM.scala 145:20:@44318.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@44319.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@44320.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@44321.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@44323.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@44322.4]
  reg  regs_37; // @[SRAM.scala 145:20:@44329.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@44330.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@44331.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@44332.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@44334.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@44333.4]
  reg  regs_38; // @[SRAM.scala 145:20:@44340.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@44341.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@44342.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@44343.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@44345.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@44344.4]
  reg  regs_39; // @[SRAM.scala 145:20:@44351.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@44352.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@44353.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@44354.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@44356.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@44355.4]
  reg  regs_40; // @[SRAM.scala 145:20:@44362.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@44363.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@44364.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@44365.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@44367.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@44366.4]
  reg  regs_41; // @[SRAM.scala 145:20:@44373.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@44374.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@44375.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@44376.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@44378.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@44377.4]
  reg  regs_42; // @[SRAM.scala 145:20:@44384.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@44385.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@44386.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@44387.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@44389.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@44388.4]
  reg  regs_43; // @[SRAM.scala 145:20:@44395.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@44396.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@44397.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@44398.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@44400.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@44399.4]
  reg  regs_44; // @[SRAM.scala 145:20:@44406.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@44407.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@44408.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@44409.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@44411.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@44410.4]
  reg  regs_45; // @[SRAM.scala 145:20:@44417.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@44418.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@44419.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@44420.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@44422.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@44421.4]
  reg  regs_46; // @[SRAM.scala 145:20:@44428.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@44429.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@44430.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@44431.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@44433.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@44432.4]
  reg  regs_47; // @[SRAM.scala 145:20:@44439.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@44440.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@44441.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@44442.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@44444.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@44443.4]
  reg  regs_48; // @[SRAM.scala 145:20:@44450.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@44451.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@44452.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@44453.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@44455.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@44454.4]
  reg  regs_49; // @[SRAM.scala 145:20:@44461.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@44462.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@44463.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@44464.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@44466.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@44465.4]
  reg  regs_50; // @[SRAM.scala 145:20:@44472.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@44473.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@44474.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@44475.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@44477.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@44476.4]
  reg  regs_51; // @[SRAM.scala 145:20:@44483.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@44484.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@44485.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@44486.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@44488.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@44487.4]
  reg  regs_52; // @[SRAM.scala 145:20:@44494.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@44495.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@44496.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@44497.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@44499.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@44498.4]
  reg  regs_53; // @[SRAM.scala 145:20:@44505.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@44506.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@44507.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@44508.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@44510.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@44509.4]
  reg  regs_54; // @[SRAM.scala 145:20:@44516.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@44517.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@44518.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@44519.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@44521.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@44520.4]
  reg  regs_55; // @[SRAM.scala 145:20:@44527.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@44528.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@44529.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@44530.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@44532.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@44531.4]
  reg  regs_56; // @[SRAM.scala 145:20:@44538.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@44539.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@44540.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@44541.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@44543.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@44542.4]
  reg  regs_57; // @[SRAM.scala 145:20:@44549.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@44550.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@44551.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@44552.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@44554.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@44553.4]
  reg  regs_58; // @[SRAM.scala 145:20:@44560.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@44561.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@44562.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@44563.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@44565.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@44564.4]
  reg  regs_59; // @[SRAM.scala 145:20:@44571.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@44572.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@44573.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@44574.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@44576.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@44575.4]
  reg  regs_60; // @[SRAM.scala 145:20:@44582.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@44583.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@44584.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@44585.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@44587.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@44586.4]
  reg  regs_61; // @[SRAM.scala 145:20:@44593.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@44594.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@44595.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@44596.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@44598.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@44597.4]
  reg  regs_62; // @[SRAM.scala 145:20:@44604.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@44605.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@44606.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@44607.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@44609.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@44608.4]
  reg  regs_63; // @[SRAM.scala 145:20:@44615.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@44616.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@44617.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@44618.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@44620.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@44619.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@44689.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@44689.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@43923.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@43924.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@43925.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43927.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@43926.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@43934.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@43935.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@43936.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43938.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@43937.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@43945.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@43946.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@43947.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43949.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@43948.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@43956.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@43957.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@43958.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43960.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@43959.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@43967.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@43968.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@43969.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43971.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@43970.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@43978.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@43979.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@43980.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43982.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@43981.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@43989.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@43990.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@43991.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43993.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@43992.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@44000.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@44001.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@44002.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44004.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@44003.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@44011.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@44012.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@44013.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44015.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@44014.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@44022.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@44023.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@44024.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44026.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@44025.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@44033.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@44034.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@44035.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44037.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@44036.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@44044.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@44045.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@44046.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44048.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@44047.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@44055.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@44056.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@44057.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44059.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@44058.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@44066.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@44067.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@44068.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44070.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@44069.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@44077.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@44078.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@44079.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44081.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@44080.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@44088.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@44089.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@44090.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44092.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@44091.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@44099.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@44100.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@44101.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44103.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@44102.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@44110.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@44111.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@44112.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44114.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@44113.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@44121.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@44122.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@44123.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44125.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@44124.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@44132.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@44133.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@44134.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44136.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@44135.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@44143.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@44144.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@44145.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44147.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@44146.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@44154.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@44155.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@44156.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44158.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@44157.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@44165.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@44166.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@44167.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44169.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@44168.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@44176.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@44177.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@44178.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44180.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@44179.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@44187.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@44188.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@44189.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44191.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@44190.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@44198.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@44199.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@44200.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44202.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@44201.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@44209.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@44210.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@44211.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44213.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@44212.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@44220.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@44221.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@44222.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44224.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@44223.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@44231.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@44232.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@44233.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44235.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@44234.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@44242.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@44243.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@44244.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44246.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@44245.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@44253.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@44254.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@44255.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44257.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@44256.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@44264.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@44265.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@44266.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44268.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@44267.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@44275.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@44276.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@44277.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44279.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@44278.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@44286.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@44287.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@44288.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44290.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@44289.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@44297.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@44298.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@44299.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44301.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@44300.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@44308.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@44309.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@44310.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44312.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@44311.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@44319.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@44320.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@44321.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44323.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@44322.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@44330.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@44331.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@44332.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44334.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@44333.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@44341.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@44342.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@44343.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44345.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@44344.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@44352.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@44353.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@44354.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44356.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@44355.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@44363.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@44364.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@44365.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44367.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@44366.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@44374.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@44375.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@44376.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44378.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@44377.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@44385.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@44386.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@44387.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44389.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@44388.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@44396.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@44397.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@44398.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44400.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@44399.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@44407.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@44408.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@44409.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44411.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@44410.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@44418.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@44419.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@44420.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44422.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@44421.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@44429.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@44430.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@44431.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44433.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@44432.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@44440.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@44441.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@44442.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44444.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@44443.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@44451.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@44452.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@44453.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44455.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@44454.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@44462.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@44463.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@44464.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44466.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@44465.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@44473.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@44474.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@44475.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44477.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@44476.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@44484.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@44485.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@44486.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44488.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@44487.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@44495.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@44496.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@44497.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44499.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@44498.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@44506.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@44507.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@44508.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44510.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@44509.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@44517.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@44518.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@44519.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44521.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@44520.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@44528.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@44529.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@44530.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44532.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@44531.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@44539.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@44540.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@44541.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44543.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@44542.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@44550.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@44551.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@44552.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44554.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@44553.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@44561.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@44562.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@44563.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44565.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@44564.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@44572.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@44573.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@44574.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44576.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@44575.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@44583.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@44584.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@44585.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44587.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@44586.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@44594.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@44595.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@44596.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44598.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@44597.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@44605.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@44606.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@44607.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44609.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@44608.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@44616.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@44617.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@44618.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44620.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@44619.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@44689.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@44689.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@44689.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@44691.2]
  input   clock, // @[:@44692.4]
  input   reset, // @[:@44693.4]
  output  io_in_ready, // @[:@44694.4]
  input   io_in_valid, // @[:@44694.4]
  input   io_in_bits, // @[:@44694.4]
  input   io_out_ready, // @[:@44694.4]
  output  io_out_valid, // @[:@44694.4]
  output  io_out_bits, // @[:@44694.4]
  input   io_banks_0_wdata_valid, // @[:@44694.4]
  input   io_banks_0_wdata_bits, // @[:@44694.4]
  input   io_banks_1_wdata_valid, // @[:@44694.4]
  input   io_banks_1_wdata_bits, // @[:@44694.4]
  input   io_banks_2_wdata_valid, // @[:@44694.4]
  input   io_banks_2_wdata_bits, // @[:@44694.4]
  input   io_banks_3_wdata_valid, // @[:@44694.4]
  input   io_banks_3_wdata_bits, // @[:@44694.4]
  input   io_banks_4_wdata_valid, // @[:@44694.4]
  input   io_banks_4_wdata_bits, // @[:@44694.4]
  input   io_banks_5_wdata_valid, // @[:@44694.4]
  input   io_banks_5_wdata_bits, // @[:@44694.4]
  input   io_banks_6_wdata_valid, // @[:@44694.4]
  input   io_banks_6_wdata_bits, // @[:@44694.4]
  input   io_banks_7_wdata_valid, // @[:@44694.4]
  input   io_banks_7_wdata_bits, // @[:@44694.4]
  input   io_banks_8_wdata_valid, // @[:@44694.4]
  input   io_banks_8_wdata_bits, // @[:@44694.4]
  input   io_banks_9_wdata_valid, // @[:@44694.4]
  input   io_banks_9_wdata_bits, // @[:@44694.4]
  input   io_banks_10_wdata_valid, // @[:@44694.4]
  input   io_banks_10_wdata_bits, // @[:@44694.4]
  input   io_banks_11_wdata_valid, // @[:@44694.4]
  input   io_banks_11_wdata_bits, // @[:@44694.4]
  input   io_banks_12_wdata_valid, // @[:@44694.4]
  input   io_banks_12_wdata_bits, // @[:@44694.4]
  input   io_banks_13_wdata_valid, // @[:@44694.4]
  input   io_banks_13_wdata_bits, // @[:@44694.4]
  input   io_banks_14_wdata_valid, // @[:@44694.4]
  input   io_banks_14_wdata_bits, // @[:@44694.4]
  input   io_banks_15_wdata_valid, // @[:@44694.4]
  input   io_banks_15_wdata_bits, // @[:@44694.4]
  input   io_banks_16_wdata_valid, // @[:@44694.4]
  input   io_banks_16_wdata_bits, // @[:@44694.4]
  input   io_banks_17_wdata_valid, // @[:@44694.4]
  input   io_banks_17_wdata_bits, // @[:@44694.4]
  input   io_banks_18_wdata_valid, // @[:@44694.4]
  input   io_banks_18_wdata_bits, // @[:@44694.4]
  input   io_banks_19_wdata_valid, // @[:@44694.4]
  input   io_banks_19_wdata_bits, // @[:@44694.4]
  input   io_banks_20_wdata_valid, // @[:@44694.4]
  input   io_banks_20_wdata_bits, // @[:@44694.4]
  input   io_banks_21_wdata_valid, // @[:@44694.4]
  input   io_banks_21_wdata_bits, // @[:@44694.4]
  input   io_banks_22_wdata_valid, // @[:@44694.4]
  input   io_banks_22_wdata_bits, // @[:@44694.4]
  input   io_banks_23_wdata_valid, // @[:@44694.4]
  input   io_banks_23_wdata_bits, // @[:@44694.4]
  input   io_banks_24_wdata_valid, // @[:@44694.4]
  input   io_banks_24_wdata_bits, // @[:@44694.4]
  input   io_banks_25_wdata_valid, // @[:@44694.4]
  input   io_banks_25_wdata_bits, // @[:@44694.4]
  input   io_banks_26_wdata_valid, // @[:@44694.4]
  input   io_banks_26_wdata_bits, // @[:@44694.4]
  input   io_banks_27_wdata_valid, // @[:@44694.4]
  input   io_banks_27_wdata_bits, // @[:@44694.4]
  input   io_banks_28_wdata_valid, // @[:@44694.4]
  input   io_banks_28_wdata_bits, // @[:@44694.4]
  input   io_banks_29_wdata_valid, // @[:@44694.4]
  input   io_banks_29_wdata_bits, // @[:@44694.4]
  input   io_banks_30_wdata_valid, // @[:@44694.4]
  input   io_banks_30_wdata_bits, // @[:@44694.4]
  input   io_banks_31_wdata_valid, // @[:@44694.4]
  input   io_banks_31_wdata_bits, // @[:@44694.4]
  input   io_banks_32_wdata_valid, // @[:@44694.4]
  input   io_banks_32_wdata_bits, // @[:@44694.4]
  input   io_banks_33_wdata_valid, // @[:@44694.4]
  input   io_banks_33_wdata_bits, // @[:@44694.4]
  input   io_banks_34_wdata_valid, // @[:@44694.4]
  input   io_banks_34_wdata_bits, // @[:@44694.4]
  input   io_banks_35_wdata_valid, // @[:@44694.4]
  input   io_banks_35_wdata_bits, // @[:@44694.4]
  input   io_banks_36_wdata_valid, // @[:@44694.4]
  input   io_banks_36_wdata_bits, // @[:@44694.4]
  input   io_banks_37_wdata_valid, // @[:@44694.4]
  input   io_banks_37_wdata_bits, // @[:@44694.4]
  input   io_banks_38_wdata_valid, // @[:@44694.4]
  input   io_banks_38_wdata_bits, // @[:@44694.4]
  input   io_banks_39_wdata_valid, // @[:@44694.4]
  input   io_banks_39_wdata_bits, // @[:@44694.4]
  input   io_banks_40_wdata_valid, // @[:@44694.4]
  input   io_banks_40_wdata_bits, // @[:@44694.4]
  input   io_banks_41_wdata_valid, // @[:@44694.4]
  input   io_banks_41_wdata_bits, // @[:@44694.4]
  input   io_banks_42_wdata_valid, // @[:@44694.4]
  input   io_banks_42_wdata_bits, // @[:@44694.4]
  input   io_banks_43_wdata_valid, // @[:@44694.4]
  input   io_banks_43_wdata_bits, // @[:@44694.4]
  input   io_banks_44_wdata_valid, // @[:@44694.4]
  input   io_banks_44_wdata_bits, // @[:@44694.4]
  input   io_banks_45_wdata_valid, // @[:@44694.4]
  input   io_banks_45_wdata_bits, // @[:@44694.4]
  input   io_banks_46_wdata_valid, // @[:@44694.4]
  input   io_banks_46_wdata_bits, // @[:@44694.4]
  input   io_banks_47_wdata_valid, // @[:@44694.4]
  input   io_banks_47_wdata_bits, // @[:@44694.4]
  input   io_banks_48_wdata_valid, // @[:@44694.4]
  input   io_banks_48_wdata_bits, // @[:@44694.4]
  input   io_banks_49_wdata_valid, // @[:@44694.4]
  input   io_banks_49_wdata_bits, // @[:@44694.4]
  input   io_banks_50_wdata_valid, // @[:@44694.4]
  input   io_banks_50_wdata_bits, // @[:@44694.4]
  input   io_banks_51_wdata_valid, // @[:@44694.4]
  input   io_banks_51_wdata_bits, // @[:@44694.4]
  input   io_banks_52_wdata_valid, // @[:@44694.4]
  input   io_banks_52_wdata_bits, // @[:@44694.4]
  input   io_banks_53_wdata_valid, // @[:@44694.4]
  input   io_banks_53_wdata_bits, // @[:@44694.4]
  input   io_banks_54_wdata_valid, // @[:@44694.4]
  input   io_banks_54_wdata_bits, // @[:@44694.4]
  input   io_banks_55_wdata_valid, // @[:@44694.4]
  input   io_banks_55_wdata_bits, // @[:@44694.4]
  input   io_banks_56_wdata_valid, // @[:@44694.4]
  input   io_banks_56_wdata_bits, // @[:@44694.4]
  input   io_banks_57_wdata_valid, // @[:@44694.4]
  input   io_banks_57_wdata_bits, // @[:@44694.4]
  input   io_banks_58_wdata_valid, // @[:@44694.4]
  input   io_banks_58_wdata_bits, // @[:@44694.4]
  input   io_banks_59_wdata_valid, // @[:@44694.4]
  input   io_banks_59_wdata_bits, // @[:@44694.4]
  input   io_banks_60_wdata_valid, // @[:@44694.4]
  input   io_banks_60_wdata_bits, // @[:@44694.4]
  input   io_banks_61_wdata_valid, // @[:@44694.4]
  input   io_banks_61_wdata_bits, // @[:@44694.4]
  input   io_banks_62_wdata_valid, // @[:@44694.4]
  input   io_banks_62_wdata_bits, // @[:@44694.4]
  input   io_banks_63_wdata_valid, // @[:@44694.4]
  input   io_banks_63_wdata_bits // @[:@44694.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@44960.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@44960.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@44960.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@44960.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@44960.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@44970.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@44970.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@44970.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@44970.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@44970.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@44985.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@44985.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@44985.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@44985.4]
  wire  writeEn; // @[FIFO.scala 30:29:@44958.4]
  wire  readEn; // @[FIFO.scala 31:29:@44959.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@44980.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@44981.4]
  wire  _T_824; // @[FIFO.scala 45:27:@44982.4]
  wire  empty; // @[FIFO.scala 45:24:@44983.4]
  wire  full; // @[FIFO.scala 46:23:@44984.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@46151.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@46152.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@44960.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@44970.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@44985.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@44958.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@44959.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@44981.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@44982.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@44983.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@44984.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@46151.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@46152.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@46158.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@46156.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@45190.4]
  assign enqCounter_clock = clock; // @[:@44961.4]
  assign enqCounter_reset = reset; // @[:@44962.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@44968.4]
  assign deqCounter_clock = clock; // @[:@44971.4]
  assign deqCounter_reset = reset; // @[:@44972.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@44978.4]
  assign FFRAM_clock = clock; // @[:@44986.4]
  assign FFRAM_reset = reset; // @[:@44987.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@45186.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@45187.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@45188.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@45189.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@45192.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@45191.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@45195.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@45194.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@45198.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@45197.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@45201.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@45200.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@45204.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@45203.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@45207.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@45206.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@45210.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@45209.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@45213.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@45212.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@45216.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@45215.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@45219.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@45218.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@45222.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@45221.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@45225.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@45224.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@45228.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@45227.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@45231.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@45230.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@45234.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@45233.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@45237.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@45236.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@45240.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@45239.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@45243.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@45242.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@45246.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@45245.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@45249.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@45248.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@45252.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@45251.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@45255.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@45254.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@45258.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@45257.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@45261.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@45260.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@45264.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@45263.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@45267.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@45266.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@45270.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@45269.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@45273.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@45272.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@45276.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@45275.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@45279.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@45278.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@45282.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@45281.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@45285.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@45284.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@45288.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@45287.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@45291.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@45290.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@45294.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@45293.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@45297.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@45296.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@45300.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@45299.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@45303.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@45302.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@45306.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@45305.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@45309.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@45308.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@45312.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@45311.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@45315.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@45314.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@45318.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@45317.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@45321.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@45320.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@45324.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@45323.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@45327.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@45326.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@45330.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@45329.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@45333.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@45332.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@45336.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@45335.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@45339.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@45338.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@45342.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@45341.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@45345.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@45344.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@45348.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@45347.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@45351.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@45350.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@45354.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@45353.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@45357.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@45356.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@45360.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@45359.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@45363.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@45362.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@45366.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@45365.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@45369.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@45368.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@45372.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@45371.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@45375.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@45374.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@45378.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@45377.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@45381.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@45380.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@46160.2]
  input         clock, // @[:@46161.4]
  input         reset, // @[:@46162.4]
  input         io_dram_cmd_ready, // @[:@46163.4]
  output        io_dram_cmd_valid, // @[:@46163.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@46163.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@46163.4]
  input         io_dram_wdata_ready, // @[:@46163.4]
  output        io_dram_wdata_valid, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@46163.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@46163.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@46163.4]
  output        io_dram_wresp_ready, // @[:@46163.4]
  input         io_dram_wresp_valid, // @[:@46163.4]
  output        io_store_cmd_ready, // @[:@46163.4]
  input         io_store_cmd_valid, // @[:@46163.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@46163.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@46163.4]
  output        io_store_data_ready, // @[:@46163.4]
  input         io_store_data_valid, // @[:@46163.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@46163.4]
  input         io_store_data_bits_wstrb, // @[:@46163.4]
  input         io_store_wresp_ready, // @[:@46163.4]
  output        io_store_wresp_valid, // @[:@46163.4]
  output        io_store_wresp_bits // @[:@46163.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@46288.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@46288.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@46288.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@46288.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@46288.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@46288.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@46288.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@46288.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@46288.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@46288.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@46694.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@46694.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@46694.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@46694.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@46694.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@46694.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@46694.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@46694.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@46694.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@46935.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@46935.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@46691.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@46288.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@46694.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@46935.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@46691.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@46688.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@46689.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@46692.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@46724.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@46725.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@46726.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@46727.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@46728.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@46729.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@46730.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@46731.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@46732.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@46733.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@46734.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@46735.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@46736.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@46737.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@46738.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@46739.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@46740.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@46870.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@46871.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@46872.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@46873.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@46874.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@46875.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@46876.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@46877.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@46878.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@46879.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@46880.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@46881.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@46882.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@46883.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@46884.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@46885.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@46886.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@46887.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@46888.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@46889.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@46890.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@46891.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@46892.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@46893.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@46894.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@46895.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@46896.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@46897.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@46898.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@46899.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@46900.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@46901.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@46902.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@46903.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@46904.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@46905.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@46906.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@46907.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@46908.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@46909.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@46910.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@46911.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@46912.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@46913.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@46914.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@46915.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@46916.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@46917.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@46918.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@46919.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@46920.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@46921.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@46922.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@46923.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@46924.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@46925.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@46926.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@46927.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@46928.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@46929.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@46930.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@46931.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@46932.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@46933.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@47202.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@46686.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@46723.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@47203.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@47204.4]
  assign cmd_clock = clock; // @[:@46289.4]
  assign cmd_reset = reset; // @[:@46290.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@46683.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@46685.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@46684.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@46687.4]
  assign wdata_clock = clock; // @[:@46695.4]
  assign wdata_reset = reset; // @[:@46696.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@46720.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@46721.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@46722.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@46934.4]
  assign wresp_clock = clock; // @[:@46936.4]
  assign wresp_reset = reset; // @[:@46937.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@47200.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@47201.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@47205.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@47271.2]
  output        io_in_ready, // @[:@47274.4]
  input         io_in_valid, // @[:@47274.4]
  input  [63:0] io_in_bits_0_addr, // @[:@47274.4]
  input  [31:0] io_in_bits_0_size, // @[:@47274.4]
  input         io_in_bits_0_isWr, // @[:@47274.4]
  input  [31:0] io_in_bits_0_tag, // @[:@47274.4]
  input         io_out_ready, // @[:@47274.4]
  output        io_out_valid, // @[:@47274.4]
  output [63:0] io_out_bits_addr, // @[:@47274.4]
  output [31:0] io_out_bits_size, // @[:@47274.4]
  output        io_out_bits_isWr, // @[:@47274.4]
  output [31:0] io_out_bits_tag // @[:@47274.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@47276.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@47276.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@47285.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@47284.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@47290.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@47289.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@47287.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@47286.4]
endmodule
module MuxPipe_1( // @[:@47292.2]
  output        io_in_ready, // @[:@47295.4]
  input         io_in_valid, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@47295.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@47295.4]
  input         io_in_bits_0_wstrb_0, // @[:@47295.4]
  input         io_in_bits_0_wstrb_1, // @[:@47295.4]
  input         io_in_bits_0_wstrb_2, // @[:@47295.4]
  input         io_in_bits_0_wstrb_3, // @[:@47295.4]
  input         io_in_bits_0_wstrb_4, // @[:@47295.4]
  input         io_in_bits_0_wstrb_5, // @[:@47295.4]
  input         io_in_bits_0_wstrb_6, // @[:@47295.4]
  input         io_in_bits_0_wstrb_7, // @[:@47295.4]
  input         io_in_bits_0_wstrb_8, // @[:@47295.4]
  input         io_in_bits_0_wstrb_9, // @[:@47295.4]
  input         io_in_bits_0_wstrb_10, // @[:@47295.4]
  input         io_in_bits_0_wstrb_11, // @[:@47295.4]
  input         io_in_bits_0_wstrb_12, // @[:@47295.4]
  input         io_in_bits_0_wstrb_13, // @[:@47295.4]
  input         io_in_bits_0_wstrb_14, // @[:@47295.4]
  input         io_in_bits_0_wstrb_15, // @[:@47295.4]
  input         io_in_bits_0_wstrb_16, // @[:@47295.4]
  input         io_in_bits_0_wstrb_17, // @[:@47295.4]
  input         io_in_bits_0_wstrb_18, // @[:@47295.4]
  input         io_in_bits_0_wstrb_19, // @[:@47295.4]
  input         io_in_bits_0_wstrb_20, // @[:@47295.4]
  input         io_in_bits_0_wstrb_21, // @[:@47295.4]
  input         io_in_bits_0_wstrb_22, // @[:@47295.4]
  input         io_in_bits_0_wstrb_23, // @[:@47295.4]
  input         io_in_bits_0_wstrb_24, // @[:@47295.4]
  input         io_in_bits_0_wstrb_25, // @[:@47295.4]
  input         io_in_bits_0_wstrb_26, // @[:@47295.4]
  input         io_in_bits_0_wstrb_27, // @[:@47295.4]
  input         io_in_bits_0_wstrb_28, // @[:@47295.4]
  input         io_in_bits_0_wstrb_29, // @[:@47295.4]
  input         io_in_bits_0_wstrb_30, // @[:@47295.4]
  input         io_in_bits_0_wstrb_31, // @[:@47295.4]
  input         io_in_bits_0_wstrb_32, // @[:@47295.4]
  input         io_in_bits_0_wstrb_33, // @[:@47295.4]
  input         io_in_bits_0_wstrb_34, // @[:@47295.4]
  input         io_in_bits_0_wstrb_35, // @[:@47295.4]
  input         io_in_bits_0_wstrb_36, // @[:@47295.4]
  input         io_in_bits_0_wstrb_37, // @[:@47295.4]
  input         io_in_bits_0_wstrb_38, // @[:@47295.4]
  input         io_in_bits_0_wstrb_39, // @[:@47295.4]
  input         io_in_bits_0_wstrb_40, // @[:@47295.4]
  input         io_in_bits_0_wstrb_41, // @[:@47295.4]
  input         io_in_bits_0_wstrb_42, // @[:@47295.4]
  input         io_in_bits_0_wstrb_43, // @[:@47295.4]
  input         io_in_bits_0_wstrb_44, // @[:@47295.4]
  input         io_in_bits_0_wstrb_45, // @[:@47295.4]
  input         io_in_bits_0_wstrb_46, // @[:@47295.4]
  input         io_in_bits_0_wstrb_47, // @[:@47295.4]
  input         io_in_bits_0_wstrb_48, // @[:@47295.4]
  input         io_in_bits_0_wstrb_49, // @[:@47295.4]
  input         io_in_bits_0_wstrb_50, // @[:@47295.4]
  input         io_in_bits_0_wstrb_51, // @[:@47295.4]
  input         io_in_bits_0_wstrb_52, // @[:@47295.4]
  input         io_in_bits_0_wstrb_53, // @[:@47295.4]
  input         io_in_bits_0_wstrb_54, // @[:@47295.4]
  input         io_in_bits_0_wstrb_55, // @[:@47295.4]
  input         io_in_bits_0_wstrb_56, // @[:@47295.4]
  input         io_in_bits_0_wstrb_57, // @[:@47295.4]
  input         io_in_bits_0_wstrb_58, // @[:@47295.4]
  input         io_in_bits_0_wstrb_59, // @[:@47295.4]
  input         io_in_bits_0_wstrb_60, // @[:@47295.4]
  input         io_in_bits_0_wstrb_61, // @[:@47295.4]
  input         io_in_bits_0_wstrb_62, // @[:@47295.4]
  input         io_in_bits_0_wstrb_63, // @[:@47295.4]
  input         io_out_ready, // @[:@47295.4]
  output        io_out_valid, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_0, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_1, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_2, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_3, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_4, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_5, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_6, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_7, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_8, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_9, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_10, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_11, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_12, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_13, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_14, // @[:@47295.4]
  output [31:0] io_out_bits_wdata_15, // @[:@47295.4]
  output        io_out_bits_wstrb_0, // @[:@47295.4]
  output        io_out_bits_wstrb_1, // @[:@47295.4]
  output        io_out_bits_wstrb_2, // @[:@47295.4]
  output        io_out_bits_wstrb_3, // @[:@47295.4]
  output        io_out_bits_wstrb_4, // @[:@47295.4]
  output        io_out_bits_wstrb_5, // @[:@47295.4]
  output        io_out_bits_wstrb_6, // @[:@47295.4]
  output        io_out_bits_wstrb_7, // @[:@47295.4]
  output        io_out_bits_wstrb_8, // @[:@47295.4]
  output        io_out_bits_wstrb_9, // @[:@47295.4]
  output        io_out_bits_wstrb_10, // @[:@47295.4]
  output        io_out_bits_wstrb_11, // @[:@47295.4]
  output        io_out_bits_wstrb_12, // @[:@47295.4]
  output        io_out_bits_wstrb_13, // @[:@47295.4]
  output        io_out_bits_wstrb_14, // @[:@47295.4]
  output        io_out_bits_wstrb_15, // @[:@47295.4]
  output        io_out_bits_wstrb_16, // @[:@47295.4]
  output        io_out_bits_wstrb_17, // @[:@47295.4]
  output        io_out_bits_wstrb_18, // @[:@47295.4]
  output        io_out_bits_wstrb_19, // @[:@47295.4]
  output        io_out_bits_wstrb_20, // @[:@47295.4]
  output        io_out_bits_wstrb_21, // @[:@47295.4]
  output        io_out_bits_wstrb_22, // @[:@47295.4]
  output        io_out_bits_wstrb_23, // @[:@47295.4]
  output        io_out_bits_wstrb_24, // @[:@47295.4]
  output        io_out_bits_wstrb_25, // @[:@47295.4]
  output        io_out_bits_wstrb_26, // @[:@47295.4]
  output        io_out_bits_wstrb_27, // @[:@47295.4]
  output        io_out_bits_wstrb_28, // @[:@47295.4]
  output        io_out_bits_wstrb_29, // @[:@47295.4]
  output        io_out_bits_wstrb_30, // @[:@47295.4]
  output        io_out_bits_wstrb_31, // @[:@47295.4]
  output        io_out_bits_wstrb_32, // @[:@47295.4]
  output        io_out_bits_wstrb_33, // @[:@47295.4]
  output        io_out_bits_wstrb_34, // @[:@47295.4]
  output        io_out_bits_wstrb_35, // @[:@47295.4]
  output        io_out_bits_wstrb_36, // @[:@47295.4]
  output        io_out_bits_wstrb_37, // @[:@47295.4]
  output        io_out_bits_wstrb_38, // @[:@47295.4]
  output        io_out_bits_wstrb_39, // @[:@47295.4]
  output        io_out_bits_wstrb_40, // @[:@47295.4]
  output        io_out_bits_wstrb_41, // @[:@47295.4]
  output        io_out_bits_wstrb_42, // @[:@47295.4]
  output        io_out_bits_wstrb_43, // @[:@47295.4]
  output        io_out_bits_wstrb_44, // @[:@47295.4]
  output        io_out_bits_wstrb_45, // @[:@47295.4]
  output        io_out_bits_wstrb_46, // @[:@47295.4]
  output        io_out_bits_wstrb_47, // @[:@47295.4]
  output        io_out_bits_wstrb_48, // @[:@47295.4]
  output        io_out_bits_wstrb_49, // @[:@47295.4]
  output        io_out_bits_wstrb_50, // @[:@47295.4]
  output        io_out_bits_wstrb_51, // @[:@47295.4]
  output        io_out_bits_wstrb_52, // @[:@47295.4]
  output        io_out_bits_wstrb_53, // @[:@47295.4]
  output        io_out_bits_wstrb_54, // @[:@47295.4]
  output        io_out_bits_wstrb_55, // @[:@47295.4]
  output        io_out_bits_wstrb_56, // @[:@47295.4]
  output        io_out_bits_wstrb_57, // @[:@47295.4]
  output        io_out_bits_wstrb_58, // @[:@47295.4]
  output        io_out_bits_wstrb_59, // @[:@47295.4]
  output        io_out_bits_wstrb_60, // @[:@47295.4]
  output        io_out_bits_wstrb_61, // @[:@47295.4]
  output        io_out_bits_wstrb_62, // @[:@47295.4]
  output        io_out_bits_wstrb_63 // @[:@47295.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@47297.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@47297.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@47382.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@47381.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@47448.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@47449.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@47450.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@47451.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@47452.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@47453.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@47454.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@47455.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@47456.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@47457.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@47458.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@47459.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@47460.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@47461.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@47462.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@47463.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@47384.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@47385.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@47386.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@47387.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@47388.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@47389.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@47390.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@47391.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@47392.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@47393.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@47394.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@47395.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@47396.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@47397.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@47398.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@47399.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@47400.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@47401.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@47402.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@47403.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@47404.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@47405.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@47406.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@47407.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@47408.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@47409.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@47410.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@47411.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@47412.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@47413.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@47414.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@47415.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@47416.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@47417.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@47418.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@47419.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@47420.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@47421.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@47422.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@47423.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@47424.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@47425.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@47426.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@47427.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@47428.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@47429.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@47430.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@47431.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@47432.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@47433.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@47434.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@47435.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@47436.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@47437.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@47438.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@47439.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@47440.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@47441.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@47442.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@47443.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@47444.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@47445.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@47446.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@47447.4]
endmodule
module ElementCounter( // @[:@47465.2]
  input         clock, // @[:@47466.4]
  input         reset, // @[:@47467.4]
  input         io_reset, // @[:@47468.4]
  input         io_enable, // @[:@47468.4]
  output [31:0] io_out // @[:@47468.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@47470.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@47471.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@47472.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@47477.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@47473.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@47471.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@47472.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@47477.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@47473.4]
  assign io_out = count; // @[Counter.scala 47:10:@47480.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@47482.2]
  input         clock, // @[:@47483.4]
  input         reset, // @[:@47484.4]
  output        io_app_0_cmd_ready, // @[:@47485.4]
  input         io_app_0_cmd_valid, // @[:@47485.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@47485.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@47485.4]
  input         io_app_0_cmd_bits_isWr, // @[:@47485.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@47485.4]
  output        io_app_0_wdata_ready, // @[:@47485.4]
  input         io_app_0_wdata_valid, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@47485.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@47485.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@47485.4]
  input         io_app_0_rresp_ready, // @[:@47485.4]
  input         io_app_0_wresp_ready, // @[:@47485.4]
  output        io_app_0_wresp_valid, // @[:@47485.4]
  input         io_dram_cmd_ready, // @[:@47485.4]
  output        io_dram_cmd_valid, // @[:@47485.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@47485.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@47485.4]
  output        io_dram_cmd_bits_isWr, // @[:@47485.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@47485.4]
  input         io_dram_wdata_ready, // @[:@47485.4]
  output        io_dram_wdata_valid, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@47485.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@47485.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@47485.4]
  output        io_dram_rresp_ready, // @[:@47485.4]
  output        io_dram_wresp_ready, // @[:@47485.4]
  input         io_dram_wresp_valid, // @[:@47485.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@47485.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47714.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47714.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@47714.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@47714.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@47714.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@47721.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@47731.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@47731.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@47731.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@47731.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@47731.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@47731.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@47731.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@47731.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@47731.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@47731.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@47731.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@47731.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@47754.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@47754.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@47757.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@47757.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@47757.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@47757.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@47757.4]
  wire  _T_346; // @[package.scala 96:25:@47726.4 package.scala 96:25:@47727.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@47728.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@47730.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@47746.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@47748.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@47751.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@47760.4]
  wire [31:0] _T_365; // @[:@47764.4 :@47765.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@47766.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@47772.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@47775.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@47776.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@47963.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@47970.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@47975.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@47979.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@47980.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@48004.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@47714.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@47721.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@47731.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@47754.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@47757.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@47726.4 package.scala 96:25:@47727.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@47728.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@47730.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@47746.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@47748.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@47751.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@47760.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@47764.4 :@47765.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@47766.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@47772.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@47775.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@47776.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@47963.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@47970.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@47975.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@47979.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@47980.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@48004.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@47977.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@47983.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@48006.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@47866.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@47865.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@47864.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@47862.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@47861.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@47949.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@47933.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@47934.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@47935.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@47936.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@47937.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@47938.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@47939.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@47940.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@47941.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@47942.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@47943.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@47944.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@47945.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@47946.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@47947.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@47948.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@47869.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@47870.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@47871.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@47872.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@47873.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@47874.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@47875.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@47876.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@47877.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@47878.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@47879.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@47880.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@47881.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@47882.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@47883.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@47884.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@47885.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@47886.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@47887.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@47888.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@47889.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@47890.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@47891.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@47892.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@47893.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@47894.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@47895.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@47896.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@47897.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@47898.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@47899.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@47900.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@47901.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@47902.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@47903.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@47904.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@47905.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@47906.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@47907.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@47908.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@47909.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@47910.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@47911.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@47912.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@47913.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@47914.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@47915.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@47916.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@47917.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@47918.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@47919.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@47920.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@47921.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@47922.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@47923.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@47924.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@47925.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@47926.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@47927.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@47928.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@47929.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@47930.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@47931.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@47932.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@48010.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@48013.4]
  assign RetimeWrapper_clock = clock; // @[:@47715.4]
  assign RetimeWrapper_reset = reset; // @[:@47716.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@47718.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@47717.4]
  assign RetimeWrapper_1_clock = clock; // @[:@47722.4]
  assign RetimeWrapper_1_reset = reset; // @[:@47723.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@47725.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@47724.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@47734.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@47740.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@47739.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@47737.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@47736.4 FringeBundles.scala 115:32:@47753.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@47867.4 StreamArbiter.scala 57:23:@47973.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@47778.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@47845.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@47846.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@47847.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@47848.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@47849.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@47850.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@47851.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@47852.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@47853.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@47854.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@47855.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@47856.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@47857.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@47858.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@47859.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@47860.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@47781.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@47782.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@47783.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@47784.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@47785.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@47786.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@47787.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@47788.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@47789.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@47790.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@47791.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@47792.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@47793.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@47794.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@47795.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@47796.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@47797.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@47798.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@47799.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@47800.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@47801.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@47802.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@47803.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@47804.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@47805.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@47806.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@47807.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@47808.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@47809.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@47810.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@47811.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@47812.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@47813.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@47814.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@47815.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@47816.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@47817.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@47818.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@47819.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@47820.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@47821.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@47822.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@47823.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@47824.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@47825.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@47826.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@47827.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@47828.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@47829.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@47830.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@47831.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@47832.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@47833.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@47834.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@47835.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@47836.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@47837.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@47838.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@47839.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@47840.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@47841.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@47842.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@47843.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@47844.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@47950.4 StreamArbiter.scala 58:25:@47974.4]
  assign elementCtr_clock = clock; // @[:@47758.4]
  assign elementCtr_reset = reset; // @[:@47759.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@47762.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@47761.4]
endmodule
module Counter_72( // @[:@48015.2]
  input         clock, // @[:@48016.4]
  input         reset, // @[:@48017.4]
  input         io_reset, // @[:@48018.4]
  input         io_enable, // @[:@48018.4]
  input  [31:0] io_stride, // @[:@48018.4]
  output [31:0] io_out, // @[:@48018.4]
  output [31:0] io_next // @[:@48018.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@48020.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@48021.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@48022.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@48027.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@48023.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@48021.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@48022.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@48027.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@48023.4]
  assign io_out = count; // @[Counter.scala 25:10:@48030.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@48031.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@48033.2]
  input         clock, // @[:@48034.4]
  input         reset, // @[:@48035.4]
  output        io_in_cmd_ready, // @[:@48036.4]
  input         io_in_cmd_valid, // @[:@48036.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@48036.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@48036.4]
  input         io_in_cmd_bits_isWr, // @[:@48036.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@48036.4]
  output        io_in_wdata_ready, // @[:@48036.4]
  input         io_in_wdata_valid, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@48036.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@48036.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@48036.4]
  input         io_in_rresp_ready, // @[:@48036.4]
  input         io_in_wresp_ready, // @[:@48036.4]
  output        io_in_wresp_valid, // @[:@48036.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@48036.4]
  input         io_out_cmd_ready, // @[:@48036.4]
  output        io_out_cmd_valid, // @[:@48036.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@48036.4]
  output [31:0] io_out_cmd_bits_size, // @[:@48036.4]
  output        io_out_cmd_bits_isWr, // @[:@48036.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@48036.4]
  input         io_out_wdata_ready, // @[:@48036.4]
  output        io_out_wdata_valid, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@48036.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@48036.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@48036.4]
  output        io_out_rresp_ready, // @[:@48036.4]
  output        io_out_wresp_ready, // @[:@48036.4]
  input         io_out_wresp_valid, // @[:@48036.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@48036.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@48150.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@48150.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@48150.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@48150.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@48150.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@48150.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@48150.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@48153.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@48154.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@48155.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@48156.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@48159.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@48159.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@48160.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@48160.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@48161.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@48164.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@48171.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@48175.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@48178.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@48181.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@48192.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@48150.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@48153.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@48154.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@48155.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@48156.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@48159.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@48159.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@48160.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@48160.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@48161.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@48164.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@48171.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@48175.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@48178.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@48181.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@48192.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@48149.4 AXIProtocol.scala 38:19:@48183.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@48142.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@48039.4 AXIProtocol.scala 46:21:@48197.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@48038.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@48148.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@48147.4 AXIProtocol.scala 29:24:@48166.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@48146.4 AXIProtocol.scala 25:24:@48158.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@48144.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@48143.4 FringeBundles.scala 115:32:@48180.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@48141.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@48125.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@48126.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@48127.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@48128.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@48129.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@48130.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@48131.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@48132.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@48133.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@48134.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@48135.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@48136.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@48137.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@48138.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@48139.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@48140.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@48061.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@48062.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@48063.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@48064.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@48065.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@48066.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@48067.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@48068.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@48069.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@48070.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@48071.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@48072.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@48073.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@48074.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@48075.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@48076.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@48077.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@48078.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@48079.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@48080.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@48081.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@48082.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@48083.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@48084.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@48085.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@48086.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@48087.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@48088.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@48089.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@48090.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@48091.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@48092.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@48093.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@48094.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@48095.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@48096.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@48097.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@48098.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@48099.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@48100.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@48101.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@48102.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@48103.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@48104.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@48105.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@48106.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@48107.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@48108.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@48109.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@48110.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@48111.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@48112.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@48113.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@48114.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@48115.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@48116.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@48117.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@48118.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@48119.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@48120.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@48121.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@48122.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@48123.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@48124.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@48059.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@48040.4 AXIProtocol.scala 47:22:@48199.4]
  assign cmdSizeCounter_clock = clock; // @[:@48151.4]
  assign cmdSizeCounter_reset = reset; // @[:@48152.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@48184.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@48185.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@48186.4]
endmodule
module AXICmdIssue( // @[:@48219.2]
  input         clock, // @[:@48220.4]
  input         reset, // @[:@48221.4]
  output        io_in_cmd_ready, // @[:@48222.4]
  input         io_in_cmd_valid, // @[:@48222.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@48222.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@48222.4]
  input         io_in_cmd_bits_isWr, // @[:@48222.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@48222.4]
  output        io_in_wdata_ready, // @[:@48222.4]
  input         io_in_wdata_valid, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@48222.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@48222.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@48222.4]
  input         io_in_rresp_ready, // @[:@48222.4]
  input         io_in_wresp_ready, // @[:@48222.4]
  output        io_in_wresp_valid, // @[:@48222.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@48222.4]
  input         io_out_cmd_ready, // @[:@48222.4]
  output        io_out_cmd_valid, // @[:@48222.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@48222.4]
  output [31:0] io_out_cmd_bits_size, // @[:@48222.4]
  output        io_out_cmd_bits_isWr, // @[:@48222.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@48222.4]
  input         io_out_wdata_ready, // @[:@48222.4]
  output        io_out_wdata_valid, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@48222.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@48222.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@48222.4]
  output        io_out_wdata_bits_wlast, // @[:@48222.4]
  output        io_out_rresp_ready, // @[:@48222.4]
  output        io_out_wresp_ready, // @[:@48222.4]
  input         io_out_wresp_valid, // @[:@48222.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@48222.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@48336.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@48336.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@48336.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@48336.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@48336.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@48336.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@48336.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@48339.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@48340.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@48341.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@48342.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@48343.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@48349.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@48350.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@48345.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@48359.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@48360.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@48336.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@48340.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@48341.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@48342.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@48343.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@48349.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@48350.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@48345.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@48359.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@48360.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@48335.4 AXIProtocol.scala 81:19:@48357.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@48328.4 AXIProtocol.scala 82:21:@48358.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@48225.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@48224.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@48334.4 AXIProtocol.scala 84:20:@48362.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@48333.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@48332.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@48330.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@48329.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@48327.4 AXIProtocol.scala 86:22:@48364.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@48311.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@48312.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@48313.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@48314.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@48315.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@48316.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@48317.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@48318.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@48319.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@48320.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@48321.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@48322.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@48323.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@48324.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@48325.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@48326.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@48247.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@48248.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@48249.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@48250.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@48251.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@48252.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@48253.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@48254.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@48255.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@48256.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@48257.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@48258.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@48259.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@48260.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@48261.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@48262.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@48263.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@48264.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@48265.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@48266.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@48267.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@48268.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@48269.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@48270.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@48271.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@48272.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@48273.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@48274.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@48275.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@48276.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@48277.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@48278.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@48279.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@48280.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@48281.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@48282.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@48283.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@48284.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@48285.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@48286.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@48287.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@48288.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@48289.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@48290.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@48291.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@48292.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@48293.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@48294.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@48295.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@48296.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@48297.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@48298.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@48299.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@48300.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@48301.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@48302.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@48303.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@48304.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@48305.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@48306.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@48307.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@48308.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@48309.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@48310.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@48246.4 AXIProtocol.scala 87:27:@48365.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@48245.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@48226.4]
  assign wdataCounter_clock = clock; // @[:@48337.4]
  assign wdataCounter_reset = reset; // @[:@48338.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@48353.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@48354.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@48355.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@48367.2]
  input         clock, // @[:@48368.4]
  input         reset, // @[:@48369.4]
  input         io_enable, // @[:@48370.4]
  output        io_app_stores_0_cmd_ready, // @[:@48370.4]
  input         io_app_stores_0_cmd_valid, // @[:@48370.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@48370.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@48370.4]
  output        io_app_stores_0_data_ready, // @[:@48370.4]
  input         io_app_stores_0_data_valid, // @[:@48370.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@48370.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@48370.4]
  input         io_app_stores_0_wresp_ready, // @[:@48370.4]
  output        io_app_stores_0_wresp_valid, // @[:@48370.4]
  output        io_app_stores_0_wresp_bits, // @[:@48370.4]
  input         io_dram_cmd_ready, // @[:@48370.4]
  output        io_dram_cmd_valid, // @[:@48370.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@48370.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@48370.4]
  output        io_dram_cmd_bits_isWr, // @[:@48370.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@48370.4]
  input         io_dram_wdata_ready, // @[:@48370.4]
  output        io_dram_wdata_valid, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@48370.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@48370.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@48370.4]
  output        io_dram_wdata_bits_wlast, // @[:@48370.4]
  output        io_dram_rresp_ready, // @[:@48370.4]
  output        io_dram_wresp_ready, // @[:@48370.4]
  input         io_dram_wresp_valid, // @[:@48370.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@48370.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@49256.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@49270.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@49498.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@49613.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@49613.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@49256.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@49270.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@49498.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@49613.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@49269.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@49265.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@49260.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@49259.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@49838.4 DRAMArbiter.scala 100:23:@49841.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@49837.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@49836.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@49834.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@49833.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@49831.4 DRAMArbiter.scala 101:25:@49843.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@49815.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@49816.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@49817.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@49818.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@49819.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@49820.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@49821.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@49822.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@49823.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@49824.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@49825.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@49826.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@49827.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@49828.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@49829.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@49830.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@49751.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@49752.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@49753.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@49754.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@49755.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@49756.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@49757.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@49758.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@49759.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@49760.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@49761.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@49762.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@49763.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@49764.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@49765.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@49766.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@49767.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@49768.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@49769.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@49770.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@49771.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@49772.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@49773.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@49774.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@49775.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@49776.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@49777.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@49778.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@49779.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@49780.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@49781.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@49782.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@49783.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@49784.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@49785.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@49786.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@49787.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@49788.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@49789.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@49790.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@49791.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@49792.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@49793.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@49794.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@49795.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@49796.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@49797.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@49798.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@49799.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@49800.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@49801.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@49802.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@49803.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@49804.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@49805.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@49806.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@49807.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@49808.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@49809.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@49810.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@49811.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@49812.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@49813.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@49814.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@49750.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@49749.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@49730.4]
  assign StreamControllerStore_clock = clock; // @[:@49257.4]
  assign StreamControllerStore_reset = reset; // @[:@49258.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@49385.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@49378.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@49275.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@49268.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@49267.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@49266.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@49264.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@49263.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@49262.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@49261.4]
  assign StreamArbiter_clock = clock; // @[:@49271.4]
  assign StreamArbiter_reset = reset; // @[:@49272.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@49496.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@49495.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@49494.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@49492.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@49491.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@49489.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@49473.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@49474.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@49475.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@49476.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@49477.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@49478.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@49479.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@49480.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@49481.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@49482.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@49483.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@49484.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@49485.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@49486.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@49487.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@49488.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@49409.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@49410.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@49411.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@49412.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@49413.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@49414.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@49415.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@49416.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@49417.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@49418.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@49419.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@49420.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@49421.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@49422.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@49423.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@49424.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@49425.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@49426.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@49427.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@49428.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@49429.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@49430.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@49431.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@49432.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@49433.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@49434.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@49435.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@49436.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@49437.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@49438.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@49439.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@49440.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@49441.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@49442.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@49443.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@49444.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@49445.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@49446.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@49447.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@49448.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@49449.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@49450.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@49451.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@49452.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@49453.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@49454.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@49455.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@49456.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@49457.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@49458.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@49459.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@49460.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@49461.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@49462.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@49463.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@49464.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@49465.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@49466.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@49467.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@49468.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@49469.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@49470.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@49471.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@49472.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@49407.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@49388.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@49612.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@49605.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@49502.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@49501.4]
  assign AXICmdSplit_clock = clock; // @[:@49499.4]
  assign AXICmdSplit_reset = reset; // @[:@49500.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@49611.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@49610.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@49609.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@49607.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@49606.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@49604.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@49588.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@49589.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@49590.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@49591.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@49592.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@49593.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@49594.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@49595.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@49596.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@49597.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@49598.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@49599.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@49600.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@49601.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@49602.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@49603.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@49524.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@49525.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@49526.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@49527.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@49528.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@49529.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@49530.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@49531.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@49532.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@49533.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@49534.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@49535.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@49536.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@49537.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@49538.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@49539.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@49540.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@49541.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@49542.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@49543.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@49544.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@49545.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@49546.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@49547.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@49548.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@49549.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@49550.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@49551.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@49552.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@49553.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@49554.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@49555.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@49556.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@49557.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@49558.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@49559.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@49560.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@49561.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@49562.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@49563.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@49564.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@49565.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@49566.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@49567.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@49568.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@49569.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@49570.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@49571.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@49572.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@49573.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@49574.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@49575.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@49576.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@49577.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@49578.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@49579.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@49580.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@49581.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@49582.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@49583.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@49584.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@49585.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@49586.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@49587.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@49522.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@49503.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@49727.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@49720.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@49617.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@49616.4]
  assign AXICmdIssue_clock = clock; // @[:@49614.4]
  assign AXICmdIssue_reset = reset; // @[:@49615.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@49726.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@49725.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@49724.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@49722.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@49721.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@49719.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@49703.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@49704.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@49705.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@49706.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@49707.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@49708.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@49709.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@49710.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@49711.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@49712.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@49713.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@49714.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@49715.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@49716.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@49717.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@49718.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@49639.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@49640.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@49641.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@49642.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@49643.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@49644.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@49645.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@49646.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@49647.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@49648.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@49649.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@49650.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@49651.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@49652.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@49653.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@49654.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@49655.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@49656.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@49657.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@49658.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@49659.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@49660.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@49661.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@49662.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@49663.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@49664.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@49665.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@49666.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@49667.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@49668.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@49669.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@49670.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@49671.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@49672.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@49673.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@49674.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@49675.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@49676.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@49677.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@49678.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@49679.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@49680.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@49681.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@49682.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@49683.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@49684.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@49685.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@49686.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@49687.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@49688.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@49689.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@49690.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@49691.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@49692.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@49693.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@49694.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@49695.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@49696.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@49697.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@49698.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@49699.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@49700.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@49701.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@49702.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@49637.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@49618.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@49839.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@49832.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@49729.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@49728.4]
endmodule
module DRAMArbiter_1( // @[:@64068.2]
  input         clock, // @[:@64069.4]
  input         reset, // @[:@64070.4]
  input         io_enable, // @[:@64071.4]
  input         io_dram_cmd_ready, // @[:@64071.4]
  output        io_dram_cmd_valid, // @[:@64071.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@64071.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@64071.4]
  output        io_dram_cmd_bits_isWr, // @[:@64071.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@64071.4]
  input         io_dram_wdata_ready, // @[:@64071.4]
  output        io_dram_wdata_valid, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@64071.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@64071.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@64071.4]
  output        io_dram_wdata_bits_wlast, // @[:@64071.4]
  output        io_dram_rresp_ready, // @[:@64071.4]
  output        io_dram_wresp_ready, // @[:@64071.4]
  input         io_dram_wresp_valid, // @[:@64071.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@64071.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@64957.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@64971.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@65199.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@65314.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@65314.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@64957.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@64971.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@65199.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@65314.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@65539.4 DRAMArbiter.scala 100:23:@65542.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@65538.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@65537.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@65535.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@65534.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@65532.4 DRAMArbiter.scala 101:25:@65544.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@65516.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@65517.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@65518.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@65519.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@65520.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@65521.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@65522.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@65523.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@65524.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@65525.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@65526.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@65527.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@65528.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@65529.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@65530.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@65531.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@65452.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@65453.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@65454.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@65455.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@65456.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@65457.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@65458.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@65459.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@65460.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@65461.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@65462.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@65463.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@65464.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@65465.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@65466.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@65467.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@65468.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@65469.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@65470.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@65471.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@65472.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@65473.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@65474.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@65475.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@65476.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@65477.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@65478.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@65479.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@65480.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@65481.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@65482.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@65483.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@65484.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@65485.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@65486.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@65487.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@65488.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@65489.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@65490.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@65491.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@65492.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@65493.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@65494.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@65495.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@65496.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@65497.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@65498.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@65499.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@65500.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@65501.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@65502.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@65503.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@65504.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@65505.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@65506.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@65507.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@65508.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@65509.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@65510.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@65511.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@65512.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@65513.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@65514.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@65515.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@65451.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@65450.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@65431.4]
  assign StreamControllerStore_clock = clock; // @[:@64958.4]
  assign StreamControllerStore_reset = reset; // @[:@64959.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@65086.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@65079.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@64976.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@64969.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@64968.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@64967.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@64965.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@64964.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@64963.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@64962.4]
  assign StreamArbiter_clock = clock; // @[:@64972.4]
  assign StreamArbiter_reset = reset; // @[:@64973.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@65197.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@65196.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@65195.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@65193.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@65192.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@65190.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@65174.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@65175.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@65176.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@65177.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@65178.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@65179.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@65180.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@65181.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@65182.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@65183.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@65184.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@65185.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@65186.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@65187.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@65188.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@65189.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@65110.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@65111.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@65112.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@65113.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@65114.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@65115.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@65116.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@65117.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@65118.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@65119.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@65120.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@65121.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@65122.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@65123.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@65124.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@65125.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@65126.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@65127.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@65128.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@65129.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@65130.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@65131.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@65132.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@65133.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@65134.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@65135.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@65136.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@65137.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@65138.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@65139.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@65140.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@65141.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@65142.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@65143.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@65144.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@65145.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@65146.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@65147.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@65148.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@65149.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@65150.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@65151.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@65152.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@65153.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@65154.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@65155.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@65156.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@65157.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@65158.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@65159.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@65160.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@65161.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@65162.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@65163.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@65164.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@65165.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@65166.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@65167.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@65168.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@65169.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@65170.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@65171.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@65172.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@65173.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@65108.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@65089.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@65313.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@65306.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@65203.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@65202.4]
  assign AXICmdSplit_clock = clock; // @[:@65200.4]
  assign AXICmdSplit_reset = reset; // @[:@65201.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@65312.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@65311.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@65310.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@65308.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@65307.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@65305.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@65289.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@65290.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@65291.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@65292.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@65293.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@65294.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@65295.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@65296.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@65297.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@65298.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@65299.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@65300.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@65301.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@65302.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@65303.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@65304.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@65225.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@65226.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@65227.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@65228.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@65229.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@65230.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@65231.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@65232.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@65233.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@65234.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@65235.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@65236.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@65237.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@65238.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@65239.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@65240.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@65241.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@65242.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@65243.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@65244.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@65245.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@65246.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@65247.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@65248.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@65249.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@65250.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@65251.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@65252.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@65253.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@65254.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@65255.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@65256.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@65257.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@65258.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@65259.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@65260.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@65261.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@65262.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@65263.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@65264.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@65265.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@65266.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@65267.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@65268.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@65269.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@65270.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@65271.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@65272.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@65273.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@65274.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@65275.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@65276.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@65277.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@65278.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@65279.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@65280.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@65281.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@65282.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@65283.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@65284.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@65285.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@65286.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@65287.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@65288.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@65223.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@65204.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@65428.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@65421.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@65318.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@65317.4]
  assign AXICmdIssue_clock = clock; // @[:@65315.4]
  assign AXICmdIssue_reset = reset; // @[:@65316.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@65427.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@65426.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@65425.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@65423.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@65422.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@65420.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@65404.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@65405.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@65406.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@65407.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@65408.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@65409.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@65410.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@65411.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@65412.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@65413.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@65414.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@65415.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@65416.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@65417.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@65418.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@65419.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@65340.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@65341.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@65342.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@65343.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@65344.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@65345.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@65346.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@65347.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@65348.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@65349.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@65350.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@65351.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@65352.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@65353.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@65354.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@65355.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@65356.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@65357.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@65358.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@65359.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@65360.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@65361.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@65362.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@65363.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@65364.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@65365.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@65366.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@65367.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@65368.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@65369.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@65370.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@65371.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@65372.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@65373.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@65374.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@65375.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@65376.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@65377.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@65378.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@65379.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@65380.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@65381.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@65382.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@65383.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@65384.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@65385.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@65386.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@65387.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@65388.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@65389.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@65390.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@65391.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@65392.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@65393.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@65394.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@65395.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@65396.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@65397.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@65398.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@65399.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@65400.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@65401.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@65402.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@65403.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@65338.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@65319.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@65540.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@65533.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@65430.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@65429.4]
endmodule
module DRAMHeap( // @[:@96176.2]
  input         io_accel_0_req_valid, // @[:@96179.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@96179.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@96179.4]
  output        io_accel_0_resp_valid, // @[:@96179.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@96179.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@96179.4]
  output        io_host_0_req_valid, // @[:@96179.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@96179.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@96179.4]
  input         io_host_0_resp_valid, // @[:@96179.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@96179.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@96179.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@96186.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@96188.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@96187.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@96183.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@96182.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@96181.4]
endmodule
module FringeFF( // @[:@96222.2]
  input         clock, // @[:@96223.4]
  input         reset, // @[:@96224.4]
  input  [63:0] io_in, // @[:@96225.4]
  input         io_reset, // @[:@96225.4]
  output [63:0] io_out, // @[:@96225.4]
  input         io_enable // @[:@96225.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@96228.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@96228.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@96228.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@96228.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@96228.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@96233.4 package.scala 96:25:@96234.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@96239.6]
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@96228.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@96233.4 package.scala 96:25:@96234.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@96239.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@96245.4]
  assign RetimeWrapper_clock = clock; // @[:@96229.4]
  assign RetimeWrapper_reset = reset; // @[:@96230.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@96232.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@96231.4]
endmodule
module MuxN( // @[:@124861.2]
  input  [63:0] io_ins_0, // @[:@124864.4]
  input  [63:0] io_ins_1, // @[:@124864.4]
  input  [63:0] io_ins_2, // @[:@124864.4]
  input  [63:0] io_ins_3, // @[:@124864.4]
  input  [63:0] io_ins_4, // @[:@124864.4]
  input  [63:0] io_ins_5, // @[:@124864.4]
  input  [63:0] io_ins_6, // @[:@124864.4]
  input  [63:0] io_ins_7, // @[:@124864.4]
  input  [63:0] io_ins_8, // @[:@124864.4]
  input  [63:0] io_ins_9, // @[:@124864.4]
  input  [63:0] io_ins_10, // @[:@124864.4]
  input  [63:0] io_ins_11, // @[:@124864.4]
  input  [63:0] io_ins_12, // @[:@124864.4]
  input  [63:0] io_ins_13, // @[:@124864.4]
  input  [63:0] io_ins_14, // @[:@124864.4]
  input  [63:0] io_ins_15, // @[:@124864.4]
  input  [63:0] io_ins_16, // @[:@124864.4]
  input  [63:0] io_ins_17, // @[:@124864.4]
  input  [63:0] io_ins_18, // @[:@124864.4]
  input  [63:0] io_ins_19, // @[:@124864.4]
  input  [63:0] io_ins_20, // @[:@124864.4]
  input  [63:0] io_ins_21, // @[:@124864.4]
  input  [63:0] io_ins_22, // @[:@124864.4]
  input  [63:0] io_ins_23, // @[:@124864.4]
  input  [63:0] io_ins_24, // @[:@124864.4]
  input  [63:0] io_ins_25, // @[:@124864.4]
  input  [63:0] io_ins_26, // @[:@124864.4]
  input  [63:0] io_ins_27, // @[:@124864.4]
  input  [63:0] io_ins_28, // @[:@124864.4]
  input  [63:0] io_ins_29, // @[:@124864.4]
  input  [63:0] io_ins_30, // @[:@124864.4]
  input  [63:0] io_ins_31, // @[:@124864.4]
  input  [63:0] io_ins_32, // @[:@124864.4]
  input  [63:0] io_ins_33, // @[:@124864.4]
  input  [63:0] io_ins_34, // @[:@124864.4]
  input  [63:0] io_ins_35, // @[:@124864.4]
  input  [63:0] io_ins_36, // @[:@124864.4]
  input  [63:0] io_ins_37, // @[:@124864.4]
  input  [63:0] io_ins_38, // @[:@124864.4]
  input  [63:0] io_ins_39, // @[:@124864.4]
  input  [63:0] io_ins_40, // @[:@124864.4]
  input  [63:0] io_ins_41, // @[:@124864.4]
  input  [63:0] io_ins_42, // @[:@124864.4]
  input  [63:0] io_ins_43, // @[:@124864.4]
  input  [63:0] io_ins_44, // @[:@124864.4]
  input  [63:0] io_ins_45, // @[:@124864.4]
  input  [63:0] io_ins_46, // @[:@124864.4]
  input  [63:0] io_ins_47, // @[:@124864.4]
  input  [63:0] io_ins_48, // @[:@124864.4]
  input  [63:0] io_ins_49, // @[:@124864.4]
  input  [63:0] io_ins_50, // @[:@124864.4]
  input  [63:0] io_ins_51, // @[:@124864.4]
  input  [63:0] io_ins_52, // @[:@124864.4]
  input  [63:0] io_ins_53, // @[:@124864.4]
  input  [63:0] io_ins_54, // @[:@124864.4]
  input  [63:0] io_ins_55, // @[:@124864.4]
  input  [63:0] io_ins_56, // @[:@124864.4]
  input  [63:0] io_ins_57, // @[:@124864.4]
  input  [63:0] io_ins_58, // @[:@124864.4]
  input  [63:0] io_ins_59, // @[:@124864.4]
  input  [63:0] io_ins_60, // @[:@124864.4]
  input  [63:0] io_ins_61, // @[:@124864.4]
  input  [63:0] io_ins_62, // @[:@124864.4]
  input  [63:0] io_ins_63, // @[:@124864.4]
  input  [63:0] io_ins_64, // @[:@124864.4]
  input  [63:0] io_ins_65, // @[:@124864.4]
  input  [63:0] io_ins_66, // @[:@124864.4]
  input  [63:0] io_ins_67, // @[:@124864.4]
  input  [63:0] io_ins_68, // @[:@124864.4]
  input  [63:0] io_ins_69, // @[:@124864.4]
  input  [63:0] io_ins_70, // @[:@124864.4]
  input  [63:0] io_ins_71, // @[:@124864.4]
  input  [63:0] io_ins_72, // @[:@124864.4]
  input  [63:0] io_ins_73, // @[:@124864.4]
  input  [63:0] io_ins_74, // @[:@124864.4]
  input  [63:0] io_ins_75, // @[:@124864.4]
  input  [63:0] io_ins_76, // @[:@124864.4]
  input  [63:0] io_ins_77, // @[:@124864.4]
  input  [63:0] io_ins_78, // @[:@124864.4]
  input  [63:0] io_ins_79, // @[:@124864.4]
  input  [63:0] io_ins_80, // @[:@124864.4]
  input  [63:0] io_ins_81, // @[:@124864.4]
  input  [63:0] io_ins_82, // @[:@124864.4]
  input  [63:0] io_ins_83, // @[:@124864.4]
  input  [63:0] io_ins_84, // @[:@124864.4]
  input  [63:0] io_ins_85, // @[:@124864.4]
  input  [63:0] io_ins_86, // @[:@124864.4]
  input  [63:0] io_ins_87, // @[:@124864.4]
  input  [63:0] io_ins_88, // @[:@124864.4]
  input  [63:0] io_ins_89, // @[:@124864.4]
  input  [63:0] io_ins_90, // @[:@124864.4]
  input  [63:0] io_ins_91, // @[:@124864.4]
  input  [63:0] io_ins_92, // @[:@124864.4]
  input  [63:0] io_ins_93, // @[:@124864.4]
  input  [63:0] io_ins_94, // @[:@124864.4]
  input  [63:0] io_ins_95, // @[:@124864.4]
  input  [63:0] io_ins_96, // @[:@124864.4]
  input  [63:0] io_ins_97, // @[:@124864.4]
  input  [63:0] io_ins_98, // @[:@124864.4]
  input  [63:0] io_ins_99, // @[:@124864.4]
  input  [63:0] io_ins_100, // @[:@124864.4]
  input  [63:0] io_ins_101, // @[:@124864.4]
  input  [63:0] io_ins_102, // @[:@124864.4]
  input  [63:0] io_ins_103, // @[:@124864.4]
  input  [63:0] io_ins_104, // @[:@124864.4]
  input  [63:0] io_ins_105, // @[:@124864.4]
  input  [63:0] io_ins_106, // @[:@124864.4]
  input  [63:0] io_ins_107, // @[:@124864.4]
  input  [63:0] io_ins_108, // @[:@124864.4]
  input  [63:0] io_ins_109, // @[:@124864.4]
  input  [63:0] io_ins_110, // @[:@124864.4]
  input  [63:0] io_ins_111, // @[:@124864.4]
  input  [63:0] io_ins_112, // @[:@124864.4]
  input  [63:0] io_ins_113, // @[:@124864.4]
  input  [63:0] io_ins_114, // @[:@124864.4]
  input  [63:0] io_ins_115, // @[:@124864.4]
  input  [63:0] io_ins_116, // @[:@124864.4]
  input  [63:0] io_ins_117, // @[:@124864.4]
  input  [63:0] io_ins_118, // @[:@124864.4]
  input  [63:0] io_ins_119, // @[:@124864.4]
  input  [63:0] io_ins_120, // @[:@124864.4]
  input  [63:0] io_ins_121, // @[:@124864.4]
  input  [63:0] io_ins_122, // @[:@124864.4]
  input  [63:0] io_ins_123, // @[:@124864.4]
  input  [63:0] io_ins_124, // @[:@124864.4]
  input  [63:0] io_ins_125, // @[:@124864.4]
  input  [63:0] io_ins_126, // @[:@124864.4]
  input  [63:0] io_ins_127, // @[:@124864.4]
  input  [63:0] io_ins_128, // @[:@124864.4]
  input  [63:0] io_ins_129, // @[:@124864.4]
  input  [63:0] io_ins_130, // @[:@124864.4]
  input  [63:0] io_ins_131, // @[:@124864.4]
  input  [63:0] io_ins_132, // @[:@124864.4]
  input  [63:0] io_ins_133, // @[:@124864.4]
  input  [63:0] io_ins_134, // @[:@124864.4]
  input  [63:0] io_ins_135, // @[:@124864.4]
  input  [63:0] io_ins_136, // @[:@124864.4]
  input  [63:0] io_ins_137, // @[:@124864.4]
  input  [63:0] io_ins_138, // @[:@124864.4]
  input  [63:0] io_ins_139, // @[:@124864.4]
  input  [63:0] io_ins_140, // @[:@124864.4]
  input  [63:0] io_ins_141, // @[:@124864.4]
  input  [63:0] io_ins_142, // @[:@124864.4]
  input  [63:0] io_ins_143, // @[:@124864.4]
  input  [63:0] io_ins_144, // @[:@124864.4]
  input  [63:0] io_ins_145, // @[:@124864.4]
  input  [63:0] io_ins_146, // @[:@124864.4]
  input  [63:0] io_ins_147, // @[:@124864.4]
  input  [63:0] io_ins_148, // @[:@124864.4]
  input  [63:0] io_ins_149, // @[:@124864.4]
  input  [63:0] io_ins_150, // @[:@124864.4]
  input  [63:0] io_ins_151, // @[:@124864.4]
  input  [63:0] io_ins_152, // @[:@124864.4]
  input  [63:0] io_ins_153, // @[:@124864.4]
  input  [63:0] io_ins_154, // @[:@124864.4]
  input  [63:0] io_ins_155, // @[:@124864.4]
  input  [63:0] io_ins_156, // @[:@124864.4]
  input  [63:0] io_ins_157, // @[:@124864.4]
  input  [63:0] io_ins_158, // @[:@124864.4]
  input  [63:0] io_ins_159, // @[:@124864.4]
  input  [63:0] io_ins_160, // @[:@124864.4]
  input  [63:0] io_ins_161, // @[:@124864.4]
  input  [63:0] io_ins_162, // @[:@124864.4]
  input  [63:0] io_ins_163, // @[:@124864.4]
  input  [63:0] io_ins_164, // @[:@124864.4]
  input  [63:0] io_ins_165, // @[:@124864.4]
  input  [63:0] io_ins_166, // @[:@124864.4]
  input  [63:0] io_ins_167, // @[:@124864.4]
  input  [63:0] io_ins_168, // @[:@124864.4]
  input  [63:0] io_ins_169, // @[:@124864.4]
  input  [63:0] io_ins_170, // @[:@124864.4]
  input  [63:0] io_ins_171, // @[:@124864.4]
  input  [63:0] io_ins_172, // @[:@124864.4]
  input  [63:0] io_ins_173, // @[:@124864.4]
  input  [63:0] io_ins_174, // @[:@124864.4]
  input  [63:0] io_ins_175, // @[:@124864.4]
  input  [63:0] io_ins_176, // @[:@124864.4]
  input  [63:0] io_ins_177, // @[:@124864.4]
  input  [63:0] io_ins_178, // @[:@124864.4]
  input  [63:0] io_ins_179, // @[:@124864.4]
  input  [63:0] io_ins_180, // @[:@124864.4]
  input  [63:0] io_ins_181, // @[:@124864.4]
  input  [63:0] io_ins_182, // @[:@124864.4]
  input  [63:0] io_ins_183, // @[:@124864.4]
  input  [63:0] io_ins_184, // @[:@124864.4]
  input  [63:0] io_ins_185, // @[:@124864.4]
  input  [63:0] io_ins_186, // @[:@124864.4]
  input  [63:0] io_ins_187, // @[:@124864.4]
  input  [63:0] io_ins_188, // @[:@124864.4]
  input  [63:0] io_ins_189, // @[:@124864.4]
  input  [63:0] io_ins_190, // @[:@124864.4]
  input  [63:0] io_ins_191, // @[:@124864.4]
  input  [63:0] io_ins_192, // @[:@124864.4]
  input  [63:0] io_ins_193, // @[:@124864.4]
  input  [63:0] io_ins_194, // @[:@124864.4]
  input  [63:0] io_ins_195, // @[:@124864.4]
  input  [63:0] io_ins_196, // @[:@124864.4]
  input  [63:0] io_ins_197, // @[:@124864.4]
  input  [63:0] io_ins_198, // @[:@124864.4]
  input  [63:0] io_ins_199, // @[:@124864.4]
  input  [63:0] io_ins_200, // @[:@124864.4]
  input  [63:0] io_ins_201, // @[:@124864.4]
  input  [63:0] io_ins_202, // @[:@124864.4]
  input  [63:0] io_ins_203, // @[:@124864.4]
  input  [63:0] io_ins_204, // @[:@124864.4]
  input  [63:0] io_ins_205, // @[:@124864.4]
  input  [63:0] io_ins_206, // @[:@124864.4]
  input  [63:0] io_ins_207, // @[:@124864.4]
  input  [63:0] io_ins_208, // @[:@124864.4]
  input  [63:0] io_ins_209, // @[:@124864.4]
  input  [63:0] io_ins_210, // @[:@124864.4]
  input  [63:0] io_ins_211, // @[:@124864.4]
  input  [63:0] io_ins_212, // @[:@124864.4]
  input  [63:0] io_ins_213, // @[:@124864.4]
  input  [63:0] io_ins_214, // @[:@124864.4]
  input  [63:0] io_ins_215, // @[:@124864.4]
  input  [63:0] io_ins_216, // @[:@124864.4]
  input  [63:0] io_ins_217, // @[:@124864.4]
  input  [63:0] io_ins_218, // @[:@124864.4]
  input  [63:0] io_ins_219, // @[:@124864.4]
  input  [63:0] io_ins_220, // @[:@124864.4]
  input  [63:0] io_ins_221, // @[:@124864.4]
  input  [63:0] io_ins_222, // @[:@124864.4]
  input  [63:0] io_ins_223, // @[:@124864.4]
  input  [63:0] io_ins_224, // @[:@124864.4]
  input  [63:0] io_ins_225, // @[:@124864.4]
  input  [63:0] io_ins_226, // @[:@124864.4]
  input  [63:0] io_ins_227, // @[:@124864.4]
  input  [63:0] io_ins_228, // @[:@124864.4]
  input  [63:0] io_ins_229, // @[:@124864.4]
  input  [63:0] io_ins_230, // @[:@124864.4]
  input  [63:0] io_ins_231, // @[:@124864.4]
  input  [63:0] io_ins_232, // @[:@124864.4]
  input  [63:0] io_ins_233, // @[:@124864.4]
  input  [63:0] io_ins_234, // @[:@124864.4]
  input  [63:0] io_ins_235, // @[:@124864.4]
  input  [63:0] io_ins_236, // @[:@124864.4]
  input  [63:0] io_ins_237, // @[:@124864.4]
  input  [63:0] io_ins_238, // @[:@124864.4]
  input  [63:0] io_ins_239, // @[:@124864.4]
  input  [63:0] io_ins_240, // @[:@124864.4]
  input  [63:0] io_ins_241, // @[:@124864.4]
  input  [63:0] io_ins_242, // @[:@124864.4]
  input  [63:0] io_ins_243, // @[:@124864.4]
  input  [63:0] io_ins_244, // @[:@124864.4]
  input  [63:0] io_ins_245, // @[:@124864.4]
  input  [63:0] io_ins_246, // @[:@124864.4]
  input  [63:0] io_ins_247, // @[:@124864.4]
  input  [63:0] io_ins_248, // @[:@124864.4]
  input  [63:0] io_ins_249, // @[:@124864.4]
  input  [63:0] io_ins_250, // @[:@124864.4]
  input  [63:0] io_ins_251, // @[:@124864.4]
  input  [63:0] io_ins_252, // @[:@124864.4]
  input  [63:0] io_ins_253, // @[:@124864.4]
  input  [63:0] io_ins_254, // @[:@124864.4]
  input  [63:0] io_ins_255, // @[:@124864.4]
  input  [63:0] io_ins_256, // @[:@124864.4]
  input  [63:0] io_ins_257, // @[:@124864.4]
  input  [63:0] io_ins_258, // @[:@124864.4]
  input  [63:0] io_ins_259, // @[:@124864.4]
  input  [63:0] io_ins_260, // @[:@124864.4]
  input  [63:0] io_ins_261, // @[:@124864.4]
  input  [63:0] io_ins_262, // @[:@124864.4]
  input  [63:0] io_ins_263, // @[:@124864.4]
  input  [63:0] io_ins_264, // @[:@124864.4]
  input  [63:0] io_ins_265, // @[:@124864.4]
  input  [63:0] io_ins_266, // @[:@124864.4]
  input  [63:0] io_ins_267, // @[:@124864.4]
  input  [63:0] io_ins_268, // @[:@124864.4]
  input  [63:0] io_ins_269, // @[:@124864.4]
  input  [63:0] io_ins_270, // @[:@124864.4]
  input  [63:0] io_ins_271, // @[:@124864.4]
  input  [63:0] io_ins_272, // @[:@124864.4]
  input  [63:0] io_ins_273, // @[:@124864.4]
  input  [63:0] io_ins_274, // @[:@124864.4]
  input  [63:0] io_ins_275, // @[:@124864.4]
  input  [63:0] io_ins_276, // @[:@124864.4]
  input  [63:0] io_ins_277, // @[:@124864.4]
  input  [63:0] io_ins_278, // @[:@124864.4]
  input  [63:0] io_ins_279, // @[:@124864.4]
  input  [63:0] io_ins_280, // @[:@124864.4]
  input  [63:0] io_ins_281, // @[:@124864.4]
  input  [63:0] io_ins_282, // @[:@124864.4]
  input  [63:0] io_ins_283, // @[:@124864.4]
  input  [63:0] io_ins_284, // @[:@124864.4]
  input  [63:0] io_ins_285, // @[:@124864.4]
  input  [63:0] io_ins_286, // @[:@124864.4]
  input  [63:0] io_ins_287, // @[:@124864.4]
  input  [63:0] io_ins_288, // @[:@124864.4]
  input  [63:0] io_ins_289, // @[:@124864.4]
  input  [63:0] io_ins_290, // @[:@124864.4]
  input  [63:0] io_ins_291, // @[:@124864.4]
  input  [63:0] io_ins_292, // @[:@124864.4]
  input  [63:0] io_ins_293, // @[:@124864.4]
  input  [63:0] io_ins_294, // @[:@124864.4]
  input  [63:0] io_ins_295, // @[:@124864.4]
  input  [63:0] io_ins_296, // @[:@124864.4]
  input  [63:0] io_ins_297, // @[:@124864.4]
  input  [63:0] io_ins_298, // @[:@124864.4]
  input  [63:0] io_ins_299, // @[:@124864.4]
  input  [63:0] io_ins_300, // @[:@124864.4]
  input  [63:0] io_ins_301, // @[:@124864.4]
  input  [63:0] io_ins_302, // @[:@124864.4]
  input  [63:0] io_ins_303, // @[:@124864.4]
  input  [63:0] io_ins_304, // @[:@124864.4]
  input  [63:0] io_ins_305, // @[:@124864.4]
  input  [63:0] io_ins_306, // @[:@124864.4]
  input  [63:0] io_ins_307, // @[:@124864.4]
  input  [63:0] io_ins_308, // @[:@124864.4]
  input  [63:0] io_ins_309, // @[:@124864.4]
  input  [63:0] io_ins_310, // @[:@124864.4]
  input  [63:0] io_ins_311, // @[:@124864.4]
  input  [63:0] io_ins_312, // @[:@124864.4]
  input  [63:0] io_ins_313, // @[:@124864.4]
  input  [63:0] io_ins_314, // @[:@124864.4]
  input  [63:0] io_ins_315, // @[:@124864.4]
  input  [63:0] io_ins_316, // @[:@124864.4]
  input  [63:0] io_ins_317, // @[:@124864.4]
  input  [63:0] io_ins_318, // @[:@124864.4]
  input  [63:0] io_ins_319, // @[:@124864.4]
  input  [63:0] io_ins_320, // @[:@124864.4]
  input  [63:0] io_ins_321, // @[:@124864.4]
  input  [63:0] io_ins_322, // @[:@124864.4]
  input  [63:0] io_ins_323, // @[:@124864.4]
  input  [63:0] io_ins_324, // @[:@124864.4]
  input  [63:0] io_ins_325, // @[:@124864.4]
  input  [63:0] io_ins_326, // @[:@124864.4]
  input  [63:0] io_ins_327, // @[:@124864.4]
  input  [63:0] io_ins_328, // @[:@124864.4]
  input  [63:0] io_ins_329, // @[:@124864.4]
  input  [63:0] io_ins_330, // @[:@124864.4]
  input  [63:0] io_ins_331, // @[:@124864.4]
  input  [63:0] io_ins_332, // @[:@124864.4]
  input  [63:0] io_ins_333, // @[:@124864.4]
  input  [63:0] io_ins_334, // @[:@124864.4]
  input  [63:0] io_ins_335, // @[:@124864.4]
  input  [63:0] io_ins_336, // @[:@124864.4]
  input  [63:0] io_ins_337, // @[:@124864.4]
  input  [63:0] io_ins_338, // @[:@124864.4]
  input  [63:0] io_ins_339, // @[:@124864.4]
  input  [63:0] io_ins_340, // @[:@124864.4]
  input  [63:0] io_ins_341, // @[:@124864.4]
  input  [63:0] io_ins_342, // @[:@124864.4]
  input  [63:0] io_ins_343, // @[:@124864.4]
  input  [63:0] io_ins_344, // @[:@124864.4]
  input  [63:0] io_ins_345, // @[:@124864.4]
  input  [63:0] io_ins_346, // @[:@124864.4]
  input  [63:0] io_ins_347, // @[:@124864.4]
  input  [63:0] io_ins_348, // @[:@124864.4]
  input  [63:0] io_ins_349, // @[:@124864.4]
  input  [63:0] io_ins_350, // @[:@124864.4]
  input  [63:0] io_ins_351, // @[:@124864.4]
  input  [63:0] io_ins_352, // @[:@124864.4]
  input  [63:0] io_ins_353, // @[:@124864.4]
  input  [63:0] io_ins_354, // @[:@124864.4]
  input  [63:0] io_ins_355, // @[:@124864.4]
  input  [63:0] io_ins_356, // @[:@124864.4]
  input  [63:0] io_ins_357, // @[:@124864.4]
  input  [63:0] io_ins_358, // @[:@124864.4]
  input  [63:0] io_ins_359, // @[:@124864.4]
  input  [63:0] io_ins_360, // @[:@124864.4]
  input  [63:0] io_ins_361, // @[:@124864.4]
  input  [63:0] io_ins_362, // @[:@124864.4]
  input  [63:0] io_ins_363, // @[:@124864.4]
  input  [63:0] io_ins_364, // @[:@124864.4]
  input  [63:0] io_ins_365, // @[:@124864.4]
  input  [63:0] io_ins_366, // @[:@124864.4]
  input  [63:0] io_ins_367, // @[:@124864.4]
  input  [63:0] io_ins_368, // @[:@124864.4]
  input  [63:0] io_ins_369, // @[:@124864.4]
  input  [63:0] io_ins_370, // @[:@124864.4]
  input  [63:0] io_ins_371, // @[:@124864.4]
  input  [63:0] io_ins_372, // @[:@124864.4]
  input  [63:0] io_ins_373, // @[:@124864.4]
  input  [63:0] io_ins_374, // @[:@124864.4]
  input  [63:0] io_ins_375, // @[:@124864.4]
  input  [63:0] io_ins_376, // @[:@124864.4]
  input  [63:0] io_ins_377, // @[:@124864.4]
  input  [63:0] io_ins_378, // @[:@124864.4]
  input  [63:0] io_ins_379, // @[:@124864.4]
  input  [63:0] io_ins_380, // @[:@124864.4]
  input  [63:0] io_ins_381, // @[:@124864.4]
  input  [63:0] io_ins_382, // @[:@124864.4]
  input  [63:0] io_ins_383, // @[:@124864.4]
  input  [63:0] io_ins_384, // @[:@124864.4]
  input  [63:0] io_ins_385, // @[:@124864.4]
  input  [63:0] io_ins_386, // @[:@124864.4]
  input  [63:0] io_ins_387, // @[:@124864.4]
  input  [63:0] io_ins_388, // @[:@124864.4]
  input  [63:0] io_ins_389, // @[:@124864.4]
  input  [63:0] io_ins_390, // @[:@124864.4]
  input  [63:0] io_ins_391, // @[:@124864.4]
  input  [63:0] io_ins_392, // @[:@124864.4]
  input  [63:0] io_ins_393, // @[:@124864.4]
  input  [63:0] io_ins_394, // @[:@124864.4]
  input  [63:0] io_ins_395, // @[:@124864.4]
  input  [63:0] io_ins_396, // @[:@124864.4]
  input  [63:0] io_ins_397, // @[:@124864.4]
  input  [63:0] io_ins_398, // @[:@124864.4]
  input  [63:0] io_ins_399, // @[:@124864.4]
  input  [63:0] io_ins_400, // @[:@124864.4]
  input  [63:0] io_ins_401, // @[:@124864.4]
  input  [63:0] io_ins_402, // @[:@124864.4]
  input  [63:0] io_ins_403, // @[:@124864.4]
  input  [63:0] io_ins_404, // @[:@124864.4]
  input  [63:0] io_ins_405, // @[:@124864.4]
  input  [63:0] io_ins_406, // @[:@124864.4]
  input  [63:0] io_ins_407, // @[:@124864.4]
  input  [63:0] io_ins_408, // @[:@124864.4]
  input  [63:0] io_ins_409, // @[:@124864.4]
  input  [63:0] io_ins_410, // @[:@124864.4]
  input  [63:0] io_ins_411, // @[:@124864.4]
  input  [63:0] io_ins_412, // @[:@124864.4]
  input  [63:0] io_ins_413, // @[:@124864.4]
  input  [63:0] io_ins_414, // @[:@124864.4]
  input  [63:0] io_ins_415, // @[:@124864.4]
  input  [63:0] io_ins_416, // @[:@124864.4]
  input  [63:0] io_ins_417, // @[:@124864.4]
  input  [63:0] io_ins_418, // @[:@124864.4]
  input  [63:0] io_ins_419, // @[:@124864.4]
  input  [63:0] io_ins_420, // @[:@124864.4]
  input  [63:0] io_ins_421, // @[:@124864.4]
  input  [63:0] io_ins_422, // @[:@124864.4]
  input  [63:0] io_ins_423, // @[:@124864.4]
  input  [63:0] io_ins_424, // @[:@124864.4]
  input  [63:0] io_ins_425, // @[:@124864.4]
  input  [63:0] io_ins_426, // @[:@124864.4]
  input  [63:0] io_ins_427, // @[:@124864.4]
  input  [63:0] io_ins_428, // @[:@124864.4]
  input  [63:0] io_ins_429, // @[:@124864.4]
  input  [63:0] io_ins_430, // @[:@124864.4]
  input  [63:0] io_ins_431, // @[:@124864.4]
  input  [63:0] io_ins_432, // @[:@124864.4]
  input  [63:0] io_ins_433, // @[:@124864.4]
  input  [63:0] io_ins_434, // @[:@124864.4]
  input  [63:0] io_ins_435, // @[:@124864.4]
  input  [63:0] io_ins_436, // @[:@124864.4]
  input  [63:0] io_ins_437, // @[:@124864.4]
  input  [63:0] io_ins_438, // @[:@124864.4]
  input  [63:0] io_ins_439, // @[:@124864.4]
  input  [63:0] io_ins_440, // @[:@124864.4]
  input  [63:0] io_ins_441, // @[:@124864.4]
  input  [63:0] io_ins_442, // @[:@124864.4]
  input  [63:0] io_ins_443, // @[:@124864.4]
  input  [63:0] io_ins_444, // @[:@124864.4]
  input  [63:0] io_ins_445, // @[:@124864.4]
  input  [63:0] io_ins_446, // @[:@124864.4]
  input  [63:0] io_ins_447, // @[:@124864.4]
  input  [63:0] io_ins_448, // @[:@124864.4]
  input  [63:0] io_ins_449, // @[:@124864.4]
  input  [63:0] io_ins_450, // @[:@124864.4]
  input  [63:0] io_ins_451, // @[:@124864.4]
  input  [63:0] io_ins_452, // @[:@124864.4]
  input  [63:0] io_ins_453, // @[:@124864.4]
  input  [63:0] io_ins_454, // @[:@124864.4]
  input  [63:0] io_ins_455, // @[:@124864.4]
  input  [63:0] io_ins_456, // @[:@124864.4]
  input  [63:0] io_ins_457, // @[:@124864.4]
  input  [63:0] io_ins_458, // @[:@124864.4]
  input  [63:0] io_ins_459, // @[:@124864.4]
  input  [63:0] io_ins_460, // @[:@124864.4]
  input  [63:0] io_ins_461, // @[:@124864.4]
  input  [63:0] io_ins_462, // @[:@124864.4]
  input  [63:0] io_ins_463, // @[:@124864.4]
  input  [63:0] io_ins_464, // @[:@124864.4]
  input  [63:0] io_ins_465, // @[:@124864.4]
  input  [63:0] io_ins_466, // @[:@124864.4]
  input  [63:0] io_ins_467, // @[:@124864.4]
  input  [63:0] io_ins_468, // @[:@124864.4]
  input  [63:0] io_ins_469, // @[:@124864.4]
  input  [63:0] io_ins_470, // @[:@124864.4]
  input  [63:0] io_ins_471, // @[:@124864.4]
  input  [63:0] io_ins_472, // @[:@124864.4]
  input  [63:0] io_ins_473, // @[:@124864.4]
  input  [63:0] io_ins_474, // @[:@124864.4]
  input  [63:0] io_ins_475, // @[:@124864.4]
  input  [63:0] io_ins_476, // @[:@124864.4]
  input  [63:0] io_ins_477, // @[:@124864.4]
  input  [63:0] io_ins_478, // @[:@124864.4]
  input  [63:0] io_ins_479, // @[:@124864.4]
  input  [63:0] io_ins_480, // @[:@124864.4]
  input  [63:0] io_ins_481, // @[:@124864.4]
  input  [63:0] io_ins_482, // @[:@124864.4]
  input  [63:0] io_ins_483, // @[:@124864.4]
  input  [63:0] io_ins_484, // @[:@124864.4]
  input  [63:0] io_ins_485, // @[:@124864.4]
  input  [63:0] io_ins_486, // @[:@124864.4]
  input  [63:0] io_ins_487, // @[:@124864.4]
  input  [63:0] io_ins_488, // @[:@124864.4]
  input  [63:0] io_ins_489, // @[:@124864.4]
  input  [63:0] io_ins_490, // @[:@124864.4]
  input  [63:0] io_ins_491, // @[:@124864.4]
  input  [63:0] io_ins_492, // @[:@124864.4]
  input  [63:0] io_ins_493, // @[:@124864.4]
  input  [63:0] io_ins_494, // @[:@124864.4]
  input  [63:0] io_ins_495, // @[:@124864.4]
  input  [63:0] io_ins_496, // @[:@124864.4]
  input  [63:0] io_ins_497, // @[:@124864.4]
  input  [63:0] io_ins_498, // @[:@124864.4]
  input  [63:0] io_ins_499, // @[:@124864.4]
  input  [63:0] io_ins_500, // @[:@124864.4]
  input  [63:0] io_ins_501, // @[:@124864.4]
  input  [63:0] io_ins_502, // @[:@124864.4]
  input  [8:0]  io_sel, // @[:@124864.4]
  output [63:0] io_out // @[:@124864.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@124866.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@124866.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@124866.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@124866.4]
endmodule
module RegFile( // @[:@124868.2]
  input         clock, // @[:@124869.4]
  input         reset, // @[:@124870.4]
  input  [31:0] io_raddr, // @[:@124871.4]
  input         io_wen, // @[:@124871.4]
  input  [31:0] io_waddr, // @[:@124871.4]
  input  [63:0] io_wdata, // @[:@124871.4]
  output [63:0] io_rdata, // @[:@124871.4]
  input         io_reset, // @[:@124871.4]
  output [63:0] io_argIns_0, // @[:@124871.4]
  output [63:0] io_argIns_1, // @[:@124871.4]
  output [63:0] io_argIns_2, // @[:@124871.4]
  output [63:0] io_argIns_3, // @[:@124871.4]
  input         io_argOuts_0_valid, // @[:@124871.4]
  input  [63:0] io_argOuts_0_bits, // @[:@124871.4]
  input         io_argOuts_1_valid, // @[:@124871.4]
  input  [63:0] io_argOuts_1_bits // @[:@124871.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@126881.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@126881.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@126881.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@126881.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@126881.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@126881.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@126893.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@126893.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@126893.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@126893.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@126893.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@126893.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@126912.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@126912.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@126924.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@126924.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@126924.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@126924.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@126924.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@126924.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@126936.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@126936.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@126950.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@126950.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@126964.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@126964.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@126978.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@126978.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@126992.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@126992.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@127006.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@127006.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@127020.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@127020.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@127034.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@127034.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@127048.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@127048.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@127062.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@127062.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@127076.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@127076.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@127090.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@127090.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@127104.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@127104.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@127118.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@127118.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@127132.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@127132.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@127146.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@127146.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@127160.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@127160.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@127174.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@127174.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@127188.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@127188.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@127202.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@127202.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@127216.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@127216.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@127230.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@127230.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@127244.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@127244.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@127258.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@127258.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@127272.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@127272.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@127286.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@127286.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@127300.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@127300.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@127314.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@127314.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@127328.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@127328.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@127342.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@127342.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@127356.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@127356.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@127370.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@127370.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@127384.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@127384.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@127398.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@127398.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@127412.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@127412.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@127426.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@127426.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@127440.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@127440.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@127454.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@127454.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@127468.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@127468.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@127482.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@127482.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@127496.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@127496.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@127510.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@127510.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@127524.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@127524.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@127538.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@127538.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@127552.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@127552.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@127566.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@127566.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@127580.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@127580.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@127594.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@127594.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@127608.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@127608.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@127622.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@127622.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@127636.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@127636.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@127650.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@127650.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@127664.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@127664.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@127678.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@127678.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@127692.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@127692.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@127706.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@127706.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@127720.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@127720.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@127734.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@127734.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@127748.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@127748.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@127762.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@127762.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@127776.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@127776.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@127790.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@127790.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@127804.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@127804.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@127818.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@127818.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@127832.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@127832.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@127846.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@127846.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@127860.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@127860.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@127874.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@127874.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@127888.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@127888.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@127902.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@127902.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@127916.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@127916.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@127930.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@127930.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@127944.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@127944.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@127958.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@127958.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@127972.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@127972.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@127986.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@127986.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@128000.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@128000.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@128014.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@128014.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@128028.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@128028.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@128042.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@128042.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@128056.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@128056.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@128070.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@128070.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@128084.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@128084.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@128098.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@128098.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@128112.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@128112.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@128126.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@128126.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@128140.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@128140.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@128154.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@128154.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@128168.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@128168.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@128182.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@128182.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@128196.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@128196.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@128210.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@128210.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@128224.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@128224.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@128238.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@128238.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@128252.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@128252.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@128266.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@128266.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@128280.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@128280.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@128294.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@128294.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@128308.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@128308.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@128322.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@128322.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@128336.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@128336.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@128350.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@128350.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@128364.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@128364.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@128378.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@128378.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@128392.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@128392.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@128406.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@128406.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@128420.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@128420.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@128434.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@128434.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@128448.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@128448.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@128462.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@128462.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@128476.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@128476.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@128490.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@128490.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@128504.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@128504.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@128518.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@128518.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@128532.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@128532.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@128546.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@128546.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@128560.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@128560.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@128574.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@128574.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@128588.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@128588.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@128602.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@128602.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@128616.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@128616.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@128630.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@128630.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@128644.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@128644.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@128658.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@128658.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@128672.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@128672.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@128686.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@128686.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@128700.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@128700.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@128714.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@128714.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@128728.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@128728.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@128742.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@128742.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@128756.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@128756.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@128770.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@128770.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@128784.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@128784.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@128798.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@128798.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@128812.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@128812.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@128826.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@128826.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@128840.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@128840.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@128854.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@128854.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@128868.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@128868.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@128882.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@128882.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@128896.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@128896.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@128910.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@128910.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@128924.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@128924.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@128938.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@128938.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@128952.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@128952.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@128966.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@128966.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@128980.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@128980.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@128994.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@128994.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@129008.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@129008.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@129022.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@129022.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@129036.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@129036.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@129050.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@129050.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@129064.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@129064.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@129078.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@129078.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@129092.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@129092.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@129106.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@129106.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@129120.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@129120.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@129134.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@129134.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@129148.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@129148.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@129162.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@129162.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@129176.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@129176.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@129190.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@129190.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@129204.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@129204.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@129218.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@129218.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@129232.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@129232.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@129246.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@129246.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@129260.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@129260.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@129274.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@129274.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@129288.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@129288.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@129302.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@129302.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@129316.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@129316.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@129330.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@129330.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@129344.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@129344.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@129358.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@129358.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@129372.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@129372.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@129386.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@129386.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@129400.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@129400.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@129414.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@129414.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@129428.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@129428.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@129442.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@129442.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@129456.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@129456.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@129470.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@129470.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@129484.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@129484.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@129498.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@129498.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@129512.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@129512.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@129526.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@129526.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@129540.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@129540.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@129554.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@129554.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@129568.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@129568.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@129582.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@129582.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@129596.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@129596.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@129610.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@129610.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@129624.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@129624.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@129638.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@129638.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@129652.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@129652.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@129666.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@129666.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@129680.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@129680.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@129694.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@129694.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@129708.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@129708.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@129722.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@129722.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@129736.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@129736.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@129750.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@129750.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@129764.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@129764.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@129778.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@129778.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@129792.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@129792.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@129806.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@129806.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@129820.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@129820.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@129834.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@129834.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@129848.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@129848.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@129862.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@129862.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@129876.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@129876.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@129890.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@129890.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@129904.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@129904.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@129918.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@129918.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@129932.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@129932.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@129946.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@129946.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@129960.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@129960.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@129974.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@129974.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@129988.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@129988.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@130002.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@130002.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@130016.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@130016.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@130030.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@130030.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@130044.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@130044.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@130058.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@130058.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@130072.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@130072.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@130086.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@130086.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@130100.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@130100.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@130114.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@130114.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@130128.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@130128.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@130142.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@130142.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@130156.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@130156.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@130170.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@130170.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@130184.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@130184.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@130198.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@130198.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@130212.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@130212.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@130226.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@130226.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@130240.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@130240.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@130254.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@130254.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@130268.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@130268.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@130282.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@130282.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@130296.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@130296.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@130310.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@130310.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@130324.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@130324.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@130338.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@130338.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@130352.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@130352.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@130366.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@130366.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@130380.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@130380.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@130394.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@130394.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@130408.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@130408.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@130422.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@130422.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@130436.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@130436.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@130450.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@130450.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@130464.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@130464.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@130478.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@130478.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@130492.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@130492.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@130506.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@130506.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@130520.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@130520.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@130534.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@130534.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@130548.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@130548.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@130562.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@130562.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@130576.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@130576.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@130590.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@130590.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@130604.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@130604.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@130618.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@130618.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@130632.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@130632.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@130646.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@130646.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@130660.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@130660.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@130674.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@130674.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@130688.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@130688.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@130702.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@130702.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@130716.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@130716.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@130730.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@130730.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@130744.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@130744.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@130758.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@130758.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@130772.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@130772.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@130786.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@130786.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@130800.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@130800.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@130814.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@130814.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@130828.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@130828.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@130842.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@130842.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@130856.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@130856.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@130870.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@130870.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@130884.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@130884.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@130898.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@130898.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@130912.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@130912.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@130926.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@130926.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@130940.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@130940.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@130954.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@130954.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@130968.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@130968.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@130982.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@130982.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@130996.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@130996.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@131010.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@131010.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@131024.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@131024.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@131038.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@131038.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@131052.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@131052.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@131066.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@131066.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@131080.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@131080.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@131094.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@131094.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@131108.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@131108.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@131122.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@131122.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@131136.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@131136.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@131150.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@131150.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@131164.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@131164.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@131178.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@131178.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@131192.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@131192.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@131206.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@131206.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@131220.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@131220.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@131234.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@131234.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@131248.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@131248.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@131262.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@131262.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@131276.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@131276.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@131290.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@131290.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@131304.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@131304.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@131318.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@131318.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@131332.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@131332.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@131346.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@131346.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@131360.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@131360.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@131374.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@131374.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@131388.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@131388.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@131402.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@131402.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@131416.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@131416.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@131430.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@131430.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@131444.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@131444.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@131458.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@131458.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@131472.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@131472.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@131486.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@131486.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@131500.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@131500.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@131514.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@131514.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@131528.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@131528.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@131542.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@131542.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@131556.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@131556.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@131570.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@131570.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@131584.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@131584.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@131598.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@131598.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@131612.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@131612.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@131626.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@131626.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@131640.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@131640.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@131654.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@131654.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@131668.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@131668.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@131682.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@131682.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@131696.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@131696.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@131710.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@131710.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@131724.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@131724.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@131738.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@131738.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@131752.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@131752.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@131766.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@131766.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@131780.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@131780.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@131794.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@131794.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@131808.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@131808.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@131822.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@131822.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@131836.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@131836.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@131850.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@131850.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@131864.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@131864.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@131878.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@131878.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@131892.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@131892.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@131906.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@131906.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@131920.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@131920.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@131934.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@131934.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@131948.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@131948.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@131962.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@131962.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@131976.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@131976.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@131990.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@131990.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@132004.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@132004.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@132018.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@132018.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@132018.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@132018.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@132018.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@132018.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@132032.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@132032.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@132032.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@132032.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@132032.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@132032.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@132046.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@132046.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@132046.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@132046.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@132046.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@132046.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@132060.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@132060.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@132060.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@132060.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@132060.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@132060.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@132074.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@132074.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@132074.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@132074.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@132074.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@132074.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@132088.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@132088.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@132088.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@132088.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@132088.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@132088.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@132102.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@132102.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@132102.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@132102.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@132102.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@132102.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@132116.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@132116.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@132116.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@132116.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@132116.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@132116.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@132130.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@132130.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@132130.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@132130.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@132130.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@132130.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@132144.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@132144.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@132144.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@132144.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@132144.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@132144.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@132158.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@132158.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@132158.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@132158.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@132158.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@132158.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@132172.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@132172.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@132172.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@132172.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@132172.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@132172.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@132186.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@132186.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@132186.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@132186.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@132186.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@132186.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@132200.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@132200.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@132200.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@132200.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@132200.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@132200.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@132214.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@132214.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@132214.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@132214.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@132214.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@132214.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@132228.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@132228.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@132228.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@132228.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@132228.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@132228.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@132242.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@132242.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@132242.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@132242.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@132242.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@132242.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@132256.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@132256.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@132256.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@132256.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@132256.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@132256.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@132270.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@132270.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@132270.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@132270.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@132270.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@132270.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@132284.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@132284.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@132284.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@132284.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@132284.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@132284.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@132298.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@132298.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@132298.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@132298.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@132298.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@132298.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@132312.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@132312.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@132312.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@132312.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@132312.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@132312.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@132326.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@132326.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@132326.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@132326.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@132326.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@132326.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@132340.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@132340.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@132340.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@132340.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@132340.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@132340.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@132354.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@132354.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@132354.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@132354.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@132354.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@132354.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@132368.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@132368.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@132368.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@132368.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@132368.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@132368.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@132382.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@132382.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@132382.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@132382.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@132382.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@132382.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@132396.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@132396.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@132396.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@132396.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@132396.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@132396.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@132410.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@132410.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@132410.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@132410.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@132410.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@132410.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@132424.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@132424.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@132424.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@132424.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@132424.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@132424.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@132438.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@132438.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@132438.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@132438.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@132438.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@132438.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@132452.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@132452.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@132452.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@132452.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@132452.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@132452.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@132466.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@132466.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@132466.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@132466.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@132466.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@132466.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@132480.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@132480.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@132480.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@132480.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@132480.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@132480.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@132494.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@132494.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@132494.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@132494.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@132494.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@132494.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@132508.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@132508.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@132508.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@132508.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@132508.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@132508.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@132522.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@132522.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@132522.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@132522.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@132522.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@132522.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@132536.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@132536.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@132536.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@132536.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@132536.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@132536.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@132550.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@132550.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@132550.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@132550.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@132550.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@132550.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@132564.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@132564.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@132564.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@132564.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@132564.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@132564.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@132578.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@132578.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@132578.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@132578.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@132578.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@132578.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@132592.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@132592.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@132592.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@132592.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@132592.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@132592.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@132606.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@132606.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@132606.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@132606.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@132606.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@132606.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@132620.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@132620.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@132620.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@132620.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@132620.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@132620.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@132634.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@132634.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@132634.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@132634.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@132634.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@132634.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@132648.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@132648.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@132648.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@132648.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@132648.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@132648.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@132662.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@132662.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@132662.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@132662.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@132662.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@132662.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@132676.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@132676.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@132676.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@132676.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@132676.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@132676.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@132690.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@132690.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@132690.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@132690.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@132690.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@132690.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@132704.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@132704.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@132704.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@132704.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@132704.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@132704.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@132718.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@132718.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@132718.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@132718.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@132718.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@132718.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@132732.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@132732.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@132732.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@132732.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@132732.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@132732.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@132746.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@132746.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@132746.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@132746.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@132746.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@132746.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@132760.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@132760.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@132760.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@132760.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@132760.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@132760.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@132774.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@132774.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@132774.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@132774.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@132774.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@132774.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@132788.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@132788.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@132788.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@132788.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@132788.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@132788.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@132802.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@132802.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@132802.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@132802.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@132802.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@132802.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@132816.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@132816.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@132816.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@132816.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@132816.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@132816.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@132830.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@132830.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@132830.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@132830.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@132830.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@132830.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@132844.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@132844.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@132844.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@132844.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@132844.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@132844.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@132858.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@132858.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@132858.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@132858.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@132858.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@132858.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@132872.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@132872.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@132872.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@132872.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@132872.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@132872.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@132886.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@132886.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@132886.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@132886.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@132886.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@132886.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@132900.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@132900.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@132900.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@132900.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@132900.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@132900.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@132914.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@132914.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@132914.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@132914.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@132914.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@132914.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@132928.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@132928.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@132928.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@132928.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@132928.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@132928.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@132942.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@132942.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@132942.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@132942.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@132942.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@132942.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@132956.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@132956.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@132956.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@132956.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@132956.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@132956.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@132970.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@132970.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@132970.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@132970.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@132970.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@132970.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@132984.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@132984.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@132984.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@132984.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@132984.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@132984.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@132998.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@132998.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@132998.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@132998.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@132998.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@132998.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@133012.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@133012.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@133012.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@133012.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@133012.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@133012.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@133026.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@133026.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@133026.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@133026.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@133026.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@133026.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@133040.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@133040.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@133040.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@133040.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@133040.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@133040.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@133054.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@133054.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@133054.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@133054.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@133054.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@133054.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@133068.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@133068.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@133068.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@133068.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@133068.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@133068.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@133082.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@133082.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@133082.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@133082.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@133082.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@133082.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@133096.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@133096.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@133096.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@133096.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@133096.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@133096.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@133110.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@133110.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@133110.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@133110.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@133110.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@133110.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@133124.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@133124.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@133124.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@133124.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@133124.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@133124.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@133138.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@133138.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@133138.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@133138.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@133138.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@133138.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@133152.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@133152.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@133152.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@133152.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@133152.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@133152.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@133166.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@133166.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@133166.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@133166.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@133166.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@133166.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@133180.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@133180.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@133180.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@133180.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@133180.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@133180.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@133194.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@133194.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@133194.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@133194.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@133194.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@133194.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@133208.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@133208.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@133208.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@133208.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@133208.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@133208.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@133222.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@133222.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@133222.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@133222.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@133222.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@133222.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@133236.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@133236.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@133236.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@133236.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@133236.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@133236.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@133250.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@133250.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@133250.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@133250.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@133250.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@133250.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@133264.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@133264.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@133264.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@133264.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@133264.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@133264.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@133278.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@133278.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@133278.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@133278.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@133278.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@133278.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@133292.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@133292.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@133292.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@133292.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@133292.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@133292.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@133306.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@133306.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@133306.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@133306.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@133306.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@133306.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@133320.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@133320.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@133320.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@133320.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@133320.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@133320.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@133334.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@133334.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@133334.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@133334.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@133334.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@133334.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@133348.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@133348.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@133348.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@133348.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@133348.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@133348.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@133362.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@133362.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@133362.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@133362.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@133362.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@133362.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@133376.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@133376.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@133376.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@133376.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@133376.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@133376.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@133390.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@133390.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@133390.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@133390.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@133390.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@133390.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@133404.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@133404.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@133404.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@133404.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@133404.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@133404.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@133418.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@133418.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@133418.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@133418.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@133418.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@133418.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@133432.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@133432.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@133432.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@133432.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@133432.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@133432.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@133446.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@133446.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@133446.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@133446.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@133446.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@133446.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@133460.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@133460.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@133460.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@133460.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@133460.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@133460.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@133474.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@133474.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@133474.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@133474.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@133474.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@133474.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@133488.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@133488.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@133488.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@133488.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@133488.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@133488.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@133502.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@133502.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@133502.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@133502.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@133502.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@133502.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@133516.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@133516.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@133516.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@133516.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@133516.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@133516.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@133530.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@133530.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@133530.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@133530.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@133530.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@133530.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@133544.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@133544.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@133544.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@133544.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@133544.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@133544.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@133558.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@133558.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@133558.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@133558.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@133558.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@133558.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@133572.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@133572.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@133572.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@133572.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@133572.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@133572.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@133586.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@133586.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@133586.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@133586.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@133586.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@133586.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@133600.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@133600.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@133600.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@133600.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@133600.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@133600.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@133614.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@133614.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@133614.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@133614.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@133614.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@133614.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@133628.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@133628.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@133628.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@133628.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@133628.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@133628.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@133642.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@133642.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@133642.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@133642.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@133642.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@133642.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@133656.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@133656.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@133656.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@133656.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@133656.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@133656.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@133670.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@133670.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@133670.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@133670.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@133670.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@133670.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@133684.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@133684.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@133684.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@133684.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@133684.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@133684.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@133698.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@133698.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@133698.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@133698.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@133698.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@133698.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@133712.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@133712.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@133712.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@133712.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@133712.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@133712.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@133726.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@133726.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@133740.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@133740.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@133740.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@133740.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@133740.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@133740.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@133754.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@133754.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@133754.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@133754.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@133754.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@133754.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@133768.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@133768.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@133768.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@133768.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@133768.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@133768.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@133782.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@133782.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@133782.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@133782.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@133782.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@133782.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@133796.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@133796.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@133796.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@133796.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@133796.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@133796.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@133810.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@133810.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@133810.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@133810.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@133810.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@133810.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@133824.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@133824.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@133824.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@133824.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@133824.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@133824.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@133838.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@133838.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@133838.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@133838.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@133838.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@133838.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@133852.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@133852.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@133852.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@133852.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@133852.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@133852.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@133866.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@133866.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@133866.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@133866.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@133866.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@133866.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@133880.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@133880.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@133880.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@133880.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@133880.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@133880.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@133894.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@133894.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@133894.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@133894.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@133894.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@133894.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@133908.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@133908.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@133908.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@133908.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@133908.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@133908.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@133922.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@133922.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@133922.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@126884.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@126896.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@126897.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@126915.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@126927.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@126939.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@126940.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@126881.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@126893.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@126912.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@126924.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@126936.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@126950.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@126964.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@126978.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@126992.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@127006.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@127020.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@127034.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@127048.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@127062.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@127076.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@127090.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@127104.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@127118.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@127132.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@127146.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@127160.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@127174.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@127188.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@127202.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@127216.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@127230.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@127244.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@127258.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@127272.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@127286.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@127300.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@127314.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@127328.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@127342.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@127356.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@127370.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@127384.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@127398.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@127412.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@127426.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@127440.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@127454.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@127468.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@127482.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@127496.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@127510.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@127524.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@127538.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@127552.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@127566.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@127580.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@127594.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@127608.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@127622.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@127636.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@127650.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@127664.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@127678.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@127692.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@127706.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@127720.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@127734.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@127748.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@127762.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@127776.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@127790.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@127804.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@127818.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@127832.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@127846.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@127860.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@127874.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@127888.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@127902.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@127916.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@127930.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@127944.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@127958.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@127972.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@127986.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@128000.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@128014.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@128028.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@128042.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@128056.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@128070.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@128084.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@128098.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@128112.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@128126.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@128140.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@128154.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@128168.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@128182.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@128196.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@128210.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@128224.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@128238.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@128252.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@128266.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@128280.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@128294.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@128308.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@128322.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@128336.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@128350.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@128364.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@128378.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@128392.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@128406.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@128420.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@128434.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@128448.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@128462.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@128476.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@128490.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@128504.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@128518.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@128532.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@128546.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@128560.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@128574.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@128588.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@128602.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@128616.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@128630.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@128644.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@128658.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@128672.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@128686.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@128700.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@128714.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@128728.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@128742.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@128756.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@128770.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@128784.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@128798.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@128812.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@128826.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@128840.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@128854.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@128868.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@128882.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@128896.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@128910.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@128924.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@128938.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@128952.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@128966.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@128980.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@128994.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@129008.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@129022.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@129036.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@129050.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@129064.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@129078.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@129092.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@129106.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@129120.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@129134.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@129148.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@129162.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@129176.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@129190.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@129204.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@129218.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@129232.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@129246.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@129260.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@129274.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@129288.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@129302.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@129316.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@129330.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@129344.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@129358.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@129372.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@129386.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@129400.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@129414.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@129428.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@129442.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@129456.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@129470.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@129484.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@129498.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@129512.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@129526.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@129540.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@129554.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@129568.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@129582.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@129596.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@129610.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@129624.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@129638.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@129652.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@129666.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@129680.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@129694.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@129708.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@129722.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@129736.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@129750.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@129764.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@129778.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@129792.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@129806.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@129820.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@129834.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@129848.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@129862.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@129876.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@129890.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@129904.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@129918.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@129932.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@129946.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@129960.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@129974.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@129988.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@130002.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@130016.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@130030.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@130044.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@130058.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@130072.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@130086.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@130100.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@130114.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@130128.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@130142.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@130156.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@130170.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@130184.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@130198.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@130212.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@130226.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@130240.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@130254.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@130268.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@130282.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@130296.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@130310.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@130324.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@130338.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@130352.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@130366.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@130380.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@130394.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@130408.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@130422.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@130436.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@130450.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@130464.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@130478.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@130492.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@130506.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@130520.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@130534.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@130548.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@130562.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@130576.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@130590.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@130604.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@130618.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@130632.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@130646.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@130660.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@130674.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@130688.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@130702.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@130716.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@130730.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@130744.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@130758.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@130772.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@130786.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@130800.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@130814.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@130828.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@130842.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@130856.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@130870.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@130884.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@130898.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@130912.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@130926.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@130940.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@130954.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@130968.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@130982.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@130996.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@131010.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@131024.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@131038.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@131052.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@131066.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@131080.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@131094.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@131108.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@131122.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@131136.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@131150.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@131164.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@131178.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@131192.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@131206.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@131220.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@131234.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@131248.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@131262.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@131276.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@131290.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@131304.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@131318.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@131332.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@131346.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@131360.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@131374.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@131388.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@131402.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@131416.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@131430.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@131444.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@131458.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@131472.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@131486.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@131500.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@131514.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@131528.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@131542.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@131556.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@131570.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@131584.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@131598.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@131612.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@131626.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@131640.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@131654.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@131668.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@131682.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@131696.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@131710.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@131724.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@131738.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@131752.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@131766.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@131780.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@131794.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@131808.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@131822.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@131836.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@131850.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@131864.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@131878.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@131892.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@131906.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@131920.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@131934.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@131948.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@131962.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@131976.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@131990.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@132004.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@132018.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@132032.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@132046.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@132060.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@132074.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@132088.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@132102.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@132116.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@132130.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@132144.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@132158.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@132172.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@132186.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@132200.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@132214.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@132228.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@132242.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@132256.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@132270.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@132284.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@132298.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@132312.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@132326.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@132340.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@132354.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@132368.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@132382.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@132396.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@132410.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@132424.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@132438.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@132452.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@132466.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@132480.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@132494.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@132508.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@132522.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@132536.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@132550.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@132564.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@132578.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@132592.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@132606.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@132620.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@132634.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@132648.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@132662.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@132676.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@132690.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@132704.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@132718.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@132732.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@132746.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@132760.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@132774.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@132788.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@132802.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@132816.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@132830.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@132844.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@132858.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@132872.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@132886.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@132900.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@132914.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@132928.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@132942.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@132956.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@132970.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@132984.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@132998.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@133012.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@133026.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@133040.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@133054.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@133068.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@133082.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@133096.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@133110.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@133124.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@133138.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@133152.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@133166.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@133180.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@133194.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@133208.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@133222.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@133236.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@133250.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@133264.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@133278.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@133292.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@133306.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@133320.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@133334.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@133348.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@133362.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@133376.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@133390.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@133404.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@133418.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@133432.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@133446.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@133460.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@133474.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@133488.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@133502.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@133516.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@133530.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@133544.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@133558.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@133572.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@133586.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@133600.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@133614.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@133628.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@133642.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@133656.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@133670.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@133684.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@133698.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@133712.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@133726.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@133740.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@133754.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@133768.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@133782.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@133796.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@133810.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@133824.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@133838.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@133852.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@133866.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@133880.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@133894.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@133908.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@133922.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@126884.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@126896.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@126897.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@126915.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@126927.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@126939.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@126940.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@134933.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@134939.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@134940.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@134941.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@134942.4]
  assign regs_0_clock = clock; // @[:@126882.4]
  assign regs_0_reset = reset; // @[:@126883.4 RegFile.scala 82:16:@126889.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@126887.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@126891.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@126886.4]
  assign regs_1_clock = clock; // @[:@126894.4]
  assign regs_1_reset = reset; // @[:@126895.4 RegFile.scala 70:16:@126907.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@126905.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@126910.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@126901.4]
  assign regs_2_clock = clock; // @[:@126913.4]
  assign regs_2_reset = reset; // @[:@126914.4 RegFile.scala 82:16:@126920.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@126918.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@126922.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@126917.4]
  assign regs_3_clock = clock; // @[:@126925.4]
  assign regs_3_reset = reset; // @[:@126926.4 RegFile.scala 82:16:@126932.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@126930.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@126934.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@126929.4]
  assign regs_4_clock = clock; // @[:@126937.4]
  assign regs_4_reset = io_reset; // @[:@126938.4 RegFile.scala 76:16:@126945.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@126944.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@126948.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@126942.4]
  assign regs_5_clock = clock; // @[:@126951.4]
  assign regs_5_reset = io_reset; // @[:@126952.4 RegFile.scala 76:16:@126959.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@126958.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@126962.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@126956.4]
  assign regs_6_clock = clock; // @[:@126965.4]
  assign regs_6_reset = io_reset; // @[:@126966.4 RegFile.scala 76:16:@126973.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@126972.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@126976.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@126970.4]
  assign regs_7_clock = clock; // @[:@126979.4]
  assign regs_7_reset = io_reset; // @[:@126980.4 RegFile.scala 76:16:@126987.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@126986.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@126990.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@126984.4]
  assign regs_8_clock = clock; // @[:@126993.4]
  assign regs_8_reset = io_reset; // @[:@126994.4 RegFile.scala 76:16:@127001.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@127000.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@127004.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@126998.4]
  assign regs_9_clock = clock; // @[:@127007.4]
  assign regs_9_reset = io_reset; // @[:@127008.4 RegFile.scala 76:16:@127015.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@127014.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@127018.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@127012.4]
  assign regs_10_clock = clock; // @[:@127021.4]
  assign regs_10_reset = io_reset; // @[:@127022.4 RegFile.scala 76:16:@127029.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@127028.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@127032.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@127026.4]
  assign regs_11_clock = clock; // @[:@127035.4]
  assign regs_11_reset = io_reset; // @[:@127036.4 RegFile.scala 76:16:@127043.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@127042.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@127046.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@127040.4]
  assign regs_12_clock = clock; // @[:@127049.4]
  assign regs_12_reset = io_reset; // @[:@127050.4 RegFile.scala 76:16:@127057.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@127056.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@127060.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@127054.4]
  assign regs_13_clock = clock; // @[:@127063.4]
  assign regs_13_reset = io_reset; // @[:@127064.4 RegFile.scala 76:16:@127071.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@127070.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@127074.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@127068.4]
  assign regs_14_clock = clock; // @[:@127077.4]
  assign regs_14_reset = io_reset; // @[:@127078.4 RegFile.scala 76:16:@127085.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@127084.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@127088.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@127082.4]
  assign regs_15_clock = clock; // @[:@127091.4]
  assign regs_15_reset = io_reset; // @[:@127092.4 RegFile.scala 76:16:@127099.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@127098.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@127102.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@127096.4]
  assign regs_16_clock = clock; // @[:@127105.4]
  assign regs_16_reset = io_reset; // @[:@127106.4 RegFile.scala 76:16:@127113.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@127112.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@127116.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@127110.4]
  assign regs_17_clock = clock; // @[:@127119.4]
  assign regs_17_reset = io_reset; // @[:@127120.4 RegFile.scala 76:16:@127127.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@127126.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@127130.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@127124.4]
  assign regs_18_clock = clock; // @[:@127133.4]
  assign regs_18_reset = io_reset; // @[:@127134.4 RegFile.scala 76:16:@127141.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@127140.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@127144.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@127138.4]
  assign regs_19_clock = clock; // @[:@127147.4]
  assign regs_19_reset = io_reset; // @[:@127148.4 RegFile.scala 76:16:@127155.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@127154.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@127158.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@127152.4]
  assign regs_20_clock = clock; // @[:@127161.4]
  assign regs_20_reset = io_reset; // @[:@127162.4 RegFile.scala 76:16:@127169.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@127168.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@127172.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@127166.4]
  assign regs_21_clock = clock; // @[:@127175.4]
  assign regs_21_reset = io_reset; // @[:@127176.4 RegFile.scala 76:16:@127183.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@127182.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@127186.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@127180.4]
  assign regs_22_clock = clock; // @[:@127189.4]
  assign regs_22_reset = io_reset; // @[:@127190.4 RegFile.scala 76:16:@127197.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@127196.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@127200.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@127194.4]
  assign regs_23_clock = clock; // @[:@127203.4]
  assign regs_23_reset = io_reset; // @[:@127204.4 RegFile.scala 76:16:@127211.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@127210.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@127214.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@127208.4]
  assign regs_24_clock = clock; // @[:@127217.4]
  assign regs_24_reset = io_reset; // @[:@127218.4 RegFile.scala 76:16:@127225.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@127224.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@127228.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@127222.4]
  assign regs_25_clock = clock; // @[:@127231.4]
  assign regs_25_reset = io_reset; // @[:@127232.4 RegFile.scala 76:16:@127239.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@127238.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@127242.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@127236.4]
  assign regs_26_clock = clock; // @[:@127245.4]
  assign regs_26_reset = io_reset; // @[:@127246.4 RegFile.scala 76:16:@127253.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@127252.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@127256.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@127250.4]
  assign regs_27_clock = clock; // @[:@127259.4]
  assign regs_27_reset = io_reset; // @[:@127260.4 RegFile.scala 76:16:@127267.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@127266.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@127270.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@127264.4]
  assign regs_28_clock = clock; // @[:@127273.4]
  assign regs_28_reset = io_reset; // @[:@127274.4 RegFile.scala 76:16:@127281.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@127280.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@127284.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@127278.4]
  assign regs_29_clock = clock; // @[:@127287.4]
  assign regs_29_reset = io_reset; // @[:@127288.4 RegFile.scala 76:16:@127295.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@127294.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@127298.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@127292.4]
  assign regs_30_clock = clock; // @[:@127301.4]
  assign regs_30_reset = io_reset; // @[:@127302.4 RegFile.scala 76:16:@127309.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@127308.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@127312.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@127306.4]
  assign regs_31_clock = clock; // @[:@127315.4]
  assign regs_31_reset = io_reset; // @[:@127316.4 RegFile.scala 76:16:@127323.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@127322.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@127326.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@127320.4]
  assign regs_32_clock = clock; // @[:@127329.4]
  assign regs_32_reset = io_reset; // @[:@127330.4 RegFile.scala 76:16:@127337.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@127336.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@127340.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@127334.4]
  assign regs_33_clock = clock; // @[:@127343.4]
  assign regs_33_reset = io_reset; // @[:@127344.4 RegFile.scala 76:16:@127351.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@127350.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@127354.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@127348.4]
  assign regs_34_clock = clock; // @[:@127357.4]
  assign regs_34_reset = io_reset; // @[:@127358.4 RegFile.scala 76:16:@127365.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@127364.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@127368.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@127362.4]
  assign regs_35_clock = clock; // @[:@127371.4]
  assign regs_35_reset = io_reset; // @[:@127372.4 RegFile.scala 76:16:@127379.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@127378.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@127382.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@127376.4]
  assign regs_36_clock = clock; // @[:@127385.4]
  assign regs_36_reset = io_reset; // @[:@127386.4 RegFile.scala 76:16:@127393.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@127392.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@127396.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@127390.4]
  assign regs_37_clock = clock; // @[:@127399.4]
  assign regs_37_reset = io_reset; // @[:@127400.4 RegFile.scala 76:16:@127407.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@127406.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@127410.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@127404.4]
  assign regs_38_clock = clock; // @[:@127413.4]
  assign regs_38_reset = io_reset; // @[:@127414.4 RegFile.scala 76:16:@127421.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@127420.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@127424.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@127418.4]
  assign regs_39_clock = clock; // @[:@127427.4]
  assign regs_39_reset = io_reset; // @[:@127428.4 RegFile.scala 76:16:@127435.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@127434.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@127438.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@127432.4]
  assign regs_40_clock = clock; // @[:@127441.4]
  assign regs_40_reset = io_reset; // @[:@127442.4 RegFile.scala 76:16:@127449.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@127448.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@127452.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@127446.4]
  assign regs_41_clock = clock; // @[:@127455.4]
  assign regs_41_reset = io_reset; // @[:@127456.4 RegFile.scala 76:16:@127463.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@127462.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@127466.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@127460.4]
  assign regs_42_clock = clock; // @[:@127469.4]
  assign regs_42_reset = io_reset; // @[:@127470.4 RegFile.scala 76:16:@127477.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@127476.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@127480.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@127474.4]
  assign regs_43_clock = clock; // @[:@127483.4]
  assign regs_43_reset = io_reset; // @[:@127484.4 RegFile.scala 76:16:@127491.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@127490.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@127494.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@127488.4]
  assign regs_44_clock = clock; // @[:@127497.4]
  assign regs_44_reset = io_reset; // @[:@127498.4 RegFile.scala 76:16:@127505.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@127504.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@127508.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@127502.4]
  assign regs_45_clock = clock; // @[:@127511.4]
  assign regs_45_reset = io_reset; // @[:@127512.4 RegFile.scala 76:16:@127519.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@127518.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@127522.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@127516.4]
  assign regs_46_clock = clock; // @[:@127525.4]
  assign regs_46_reset = io_reset; // @[:@127526.4 RegFile.scala 76:16:@127533.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@127532.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@127536.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@127530.4]
  assign regs_47_clock = clock; // @[:@127539.4]
  assign regs_47_reset = io_reset; // @[:@127540.4 RegFile.scala 76:16:@127547.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@127546.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@127550.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@127544.4]
  assign regs_48_clock = clock; // @[:@127553.4]
  assign regs_48_reset = io_reset; // @[:@127554.4 RegFile.scala 76:16:@127561.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@127560.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@127564.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@127558.4]
  assign regs_49_clock = clock; // @[:@127567.4]
  assign regs_49_reset = io_reset; // @[:@127568.4 RegFile.scala 76:16:@127575.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@127574.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@127578.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@127572.4]
  assign regs_50_clock = clock; // @[:@127581.4]
  assign regs_50_reset = io_reset; // @[:@127582.4 RegFile.scala 76:16:@127589.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@127588.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@127592.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@127586.4]
  assign regs_51_clock = clock; // @[:@127595.4]
  assign regs_51_reset = io_reset; // @[:@127596.4 RegFile.scala 76:16:@127603.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@127602.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@127606.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@127600.4]
  assign regs_52_clock = clock; // @[:@127609.4]
  assign regs_52_reset = io_reset; // @[:@127610.4 RegFile.scala 76:16:@127617.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@127616.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@127620.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@127614.4]
  assign regs_53_clock = clock; // @[:@127623.4]
  assign regs_53_reset = io_reset; // @[:@127624.4 RegFile.scala 76:16:@127631.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@127630.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@127634.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@127628.4]
  assign regs_54_clock = clock; // @[:@127637.4]
  assign regs_54_reset = io_reset; // @[:@127638.4 RegFile.scala 76:16:@127645.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@127644.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@127648.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@127642.4]
  assign regs_55_clock = clock; // @[:@127651.4]
  assign regs_55_reset = io_reset; // @[:@127652.4 RegFile.scala 76:16:@127659.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@127658.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@127662.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@127656.4]
  assign regs_56_clock = clock; // @[:@127665.4]
  assign regs_56_reset = io_reset; // @[:@127666.4 RegFile.scala 76:16:@127673.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@127672.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@127676.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@127670.4]
  assign regs_57_clock = clock; // @[:@127679.4]
  assign regs_57_reset = io_reset; // @[:@127680.4 RegFile.scala 76:16:@127687.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@127686.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@127690.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@127684.4]
  assign regs_58_clock = clock; // @[:@127693.4]
  assign regs_58_reset = io_reset; // @[:@127694.4 RegFile.scala 76:16:@127701.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@127700.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@127704.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@127698.4]
  assign regs_59_clock = clock; // @[:@127707.4]
  assign regs_59_reset = io_reset; // @[:@127708.4 RegFile.scala 76:16:@127715.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@127714.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@127718.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@127712.4]
  assign regs_60_clock = clock; // @[:@127721.4]
  assign regs_60_reset = io_reset; // @[:@127722.4 RegFile.scala 76:16:@127729.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@127728.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@127732.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@127726.4]
  assign regs_61_clock = clock; // @[:@127735.4]
  assign regs_61_reset = io_reset; // @[:@127736.4 RegFile.scala 76:16:@127743.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@127742.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@127746.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@127740.4]
  assign regs_62_clock = clock; // @[:@127749.4]
  assign regs_62_reset = io_reset; // @[:@127750.4 RegFile.scala 76:16:@127757.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@127756.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@127760.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@127754.4]
  assign regs_63_clock = clock; // @[:@127763.4]
  assign regs_63_reset = io_reset; // @[:@127764.4 RegFile.scala 76:16:@127771.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@127770.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@127774.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@127768.4]
  assign regs_64_clock = clock; // @[:@127777.4]
  assign regs_64_reset = io_reset; // @[:@127778.4 RegFile.scala 76:16:@127785.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@127784.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@127788.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@127782.4]
  assign regs_65_clock = clock; // @[:@127791.4]
  assign regs_65_reset = io_reset; // @[:@127792.4 RegFile.scala 76:16:@127799.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@127798.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@127802.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@127796.4]
  assign regs_66_clock = clock; // @[:@127805.4]
  assign regs_66_reset = io_reset; // @[:@127806.4 RegFile.scala 76:16:@127813.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@127812.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@127816.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@127810.4]
  assign regs_67_clock = clock; // @[:@127819.4]
  assign regs_67_reset = io_reset; // @[:@127820.4 RegFile.scala 76:16:@127827.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@127826.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@127830.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@127824.4]
  assign regs_68_clock = clock; // @[:@127833.4]
  assign regs_68_reset = io_reset; // @[:@127834.4 RegFile.scala 76:16:@127841.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@127840.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@127844.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@127838.4]
  assign regs_69_clock = clock; // @[:@127847.4]
  assign regs_69_reset = io_reset; // @[:@127848.4 RegFile.scala 76:16:@127855.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@127854.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@127858.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@127852.4]
  assign regs_70_clock = clock; // @[:@127861.4]
  assign regs_70_reset = io_reset; // @[:@127862.4 RegFile.scala 76:16:@127869.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@127868.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@127872.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@127866.4]
  assign regs_71_clock = clock; // @[:@127875.4]
  assign regs_71_reset = io_reset; // @[:@127876.4 RegFile.scala 76:16:@127883.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@127882.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@127886.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@127880.4]
  assign regs_72_clock = clock; // @[:@127889.4]
  assign regs_72_reset = io_reset; // @[:@127890.4 RegFile.scala 76:16:@127897.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@127896.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@127900.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@127894.4]
  assign regs_73_clock = clock; // @[:@127903.4]
  assign regs_73_reset = io_reset; // @[:@127904.4 RegFile.scala 76:16:@127911.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@127910.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@127914.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@127908.4]
  assign regs_74_clock = clock; // @[:@127917.4]
  assign regs_74_reset = io_reset; // @[:@127918.4 RegFile.scala 76:16:@127925.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@127924.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@127928.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@127922.4]
  assign regs_75_clock = clock; // @[:@127931.4]
  assign regs_75_reset = io_reset; // @[:@127932.4 RegFile.scala 76:16:@127939.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@127938.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@127942.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@127936.4]
  assign regs_76_clock = clock; // @[:@127945.4]
  assign regs_76_reset = io_reset; // @[:@127946.4 RegFile.scala 76:16:@127953.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@127952.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@127956.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@127950.4]
  assign regs_77_clock = clock; // @[:@127959.4]
  assign regs_77_reset = io_reset; // @[:@127960.4 RegFile.scala 76:16:@127967.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@127966.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@127970.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@127964.4]
  assign regs_78_clock = clock; // @[:@127973.4]
  assign regs_78_reset = io_reset; // @[:@127974.4 RegFile.scala 76:16:@127981.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@127980.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@127984.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@127978.4]
  assign regs_79_clock = clock; // @[:@127987.4]
  assign regs_79_reset = io_reset; // @[:@127988.4 RegFile.scala 76:16:@127995.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@127994.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@127998.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@127992.4]
  assign regs_80_clock = clock; // @[:@128001.4]
  assign regs_80_reset = io_reset; // @[:@128002.4 RegFile.scala 76:16:@128009.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@128008.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@128012.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@128006.4]
  assign regs_81_clock = clock; // @[:@128015.4]
  assign regs_81_reset = io_reset; // @[:@128016.4 RegFile.scala 76:16:@128023.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@128022.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@128026.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@128020.4]
  assign regs_82_clock = clock; // @[:@128029.4]
  assign regs_82_reset = io_reset; // @[:@128030.4 RegFile.scala 76:16:@128037.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@128036.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@128040.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@128034.4]
  assign regs_83_clock = clock; // @[:@128043.4]
  assign regs_83_reset = io_reset; // @[:@128044.4 RegFile.scala 76:16:@128051.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@128050.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@128054.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@128048.4]
  assign regs_84_clock = clock; // @[:@128057.4]
  assign regs_84_reset = io_reset; // @[:@128058.4 RegFile.scala 76:16:@128065.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@128064.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@128068.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@128062.4]
  assign regs_85_clock = clock; // @[:@128071.4]
  assign regs_85_reset = io_reset; // @[:@128072.4 RegFile.scala 76:16:@128079.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@128078.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@128082.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@128076.4]
  assign regs_86_clock = clock; // @[:@128085.4]
  assign regs_86_reset = io_reset; // @[:@128086.4 RegFile.scala 76:16:@128093.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@128092.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@128096.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@128090.4]
  assign regs_87_clock = clock; // @[:@128099.4]
  assign regs_87_reset = io_reset; // @[:@128100.4 RegFile.scala 76:16:@128107.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@128106.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@128110.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@128104.4]
  assign regs_88_clock = clock; // @[:@128113.4]
  assign regs_88_reset = io_reset; // @[:@128114.4 RegFile.scala 76:16:@128121.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@128120.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@128124.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@128118.4]
  assign regs_89_clock = clock; // @[:@128127.4]
  assign regs_89_reset = io_reset; // @[:@128128.4 RegFile.scala 76:16:@128135.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@128134.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@128138.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@128132.4]
  assign regs_90_clock = clock; // @[:@128141.4]
  assign regs_90_reset = io_reset; // @[:@128142.4 RegFile.scala 76:16:@128149.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@128148.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@128152.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@128146.4]
  assign regs_91_clock = clock; // @[:@128155.4]
  assign regs_91_reset = io_reset; // @[:@128156.4 RegFile.scala 76:16:@128163.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@128162.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@128166.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@128160.4]
  assign regs_92_clock = clock; // @[:@128169.4]
  assign regs_92_reset = io_reset; // @[:@128170.4 RegFile.scala 76:16:@128177.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@128176.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@128180.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@128174.4]
  assign regs_93_clock = clock; // @[:@128183.4]
  assign regs_93_reset = io_reset; // @[:@128184.4 RegFile.scala 76:16:@128191.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@128190.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@128194.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@128188.4]
  assign regs_94_clock = clock; // @[:@128197.4]
  assign regs_94_reset = io_reset; // @[:@128198.4 RegFile.scala 76:16:@128205.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@128204.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@128208.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@128202.4]
  assign regs_95_clock = clock; // @[:@128211.4]
  assign regs_95_reset = io_reset; // @[:@128212.4 RegFile.scala 76:16:@128219.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@128218.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@128222.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@128216.4]
  assign regs_96_clock = clock; // @[:@128225.4]
  assign regs_96_reset = io_reset; // @[:@128226.4 RegFile.scala 76:16:@128233.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@128232.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@128236.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@128230.4]
  assign regs_97_clock = clock; // @[:@128239.4]
  assign regs_97_reset = io_reset; // @[:@128240.4 RegFile.scala 76:16:@128247.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@128246.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@128250.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@128244.4]
  assign regs_98_clock = clock; // @[:@128253.4]
  assign regs_98_reset = io_reset; // @[:@128254.4 RegFile.scala 76:16:@128261.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@128260.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@128264.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@128258.4]
  assign regs_99_clock = clock; // @[:@128267.4]
  assign regs_99_reset = io_reset; // @[:@128268.4 RegFile.scala 76:16:@128275.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@128274.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@128278.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@128272.4]
  assign regs_100_clock = clock; // @[:@128281.4]
  assign regs_100_reset = io_reset; // @[:@128282.4 RegFile.scala 76:16:@128289.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@128288.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@128292.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@128286.4]
  assign regs_101_clock = clock; // @[:@128295.4]
  assign regs_101_reset = io_reset; // @[:@128296.4 RegFile.scala 76:16:@128303.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@128302.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@128306.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@128300.4]
  assign regs_102_clock = clock; // @[:@128309.4]
  assign regs_102_reset = io_reset; // @[:@128310.4 RegFile.scala 76:16:@128317.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@128316.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@128320.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@128314.4]
  assign regs_103_clock = clock; // @[:@128323.4]
  assign regs_103_reset = io_reset; // @[:@128324.4 RegFile.scala 76:16:@128331.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@128330.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@128334.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@128328.4]
  assign regs_104_clock = clock; // @[:@128337.4]
  assign regs_104_reset = io_reset; // @[:@128338.4 RegFile.scala 76:16:@128345.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@128344.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@128348.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@128342.4]
  assign regs_105_clock = clock; // @[:@128351.4]
  assign regs_105_reset = io_reset; // @[:@128352.4 RegFile.scala 76:16:@128359.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@128358.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@128362.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@128356.4]
  assign regs_106_clock = clock; // @[:@128365.4]
  assign regs_106_reset = io_reset; // @[:@128366.4 RegFile.scala 76:16:@128373.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@128372.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@128376.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@128370.4]
  assign regs_107_clock = clock; // @[:@128379.4]
  assign regs_107_reset = io_reset; // @[:@128380.4 RegFile.scala 76:16:@128387.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@128386.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@128390.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@128384.4]
  assign regs_108_clock = clock; // @[:@128393.4]
  assign regs_108_reset = io_reset; // @[:@128394.4 RegFile.scala 76:16:@128401.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@128400.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@128404.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@128398.4]
  assign regs_109_clock = clock; // @[:@128407.4]
  assign regs_109_reset = io_reset; // @[:@128408.4 RegFile.scala 76:16:@128415.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@128414.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@128418.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@128412.4]
  assign regs_110_clock = clock; // @[:@128421.4]
  assign regs_110_reset = io_reset; // @[:@128422.4 RegFile.scala 76:16:@128429.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@128428.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@128432.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@128426.4]
  assign regs_111_clock = clock; // @[:@128435.4]
  assign regs_111_reset = io_reset; // @[:@128436.4 RegFile.scala 76:16:@128443.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@128442.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@128446.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@128440.4]
  assign regs_112_clock = clock; // @[:@128449.4]
  assign regs_112_reset = io_reset; // @[:@128450.4 RegFile.scala 76:16:@128457.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@128456.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@128460.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@128454.4]
  assign regs_113_clock = clock; // @[:@128463.4]
  assign regs_113_reset = io_reset; // @[:@128464.4 RegFile.scala 76:16:@128471.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@128470.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@128474.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@128468.4]
  assign regs_114_clock = clock; // @[:@128477.4]
  assign regs_114_reset = io_reset; // @[:@128478.4 RegFile.scala 76:16:@128485.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@128484.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@128488.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@128482.4]
  assign regs_115_clock = clock; // @[:@128491.4]
  assign regs_115_reset = io_reset; // @[:@128492.4 RegFile.scala 76:16:@128499.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@128498.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@128502.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@128496.4]
  assign regs_116_clock = clock; // @[:@128505.4]
  assign regs_116_reset = io_reset; // @[:@128506.4 RegFile.scala 76:16:@128513.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@128512.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@128516.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@128510.4]
  assign regs_117_clock = clock; // @[:@128519.4]
  assign regs_117_reset = io_reset; // @[:@128520.4 RegFile.scala 76:16:@128527.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@128526.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@128530.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@128524.4]
  assign regs_118_clock = clock; // @[:@128533.4]
  assign regs_118_reset = io_reset; // @[:@128534.4 RegFile.scala 76:16:@128541.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@128540.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@128544.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@128538.4]
  assign regs_119_clock = clock; // @[:@128547.4]
  assign regs_119_reset = io_reset; // @[:@128548.4 RegFile.scala 76:16:@128555.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@128554.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@128558.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@128552.4]
  assign regs_120_clock = clock; // @[:@128561.4]
  assign regs_120_reset = io_reset; // @[:@128562.4 RegFile.scala 76:16:@128569.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@128568.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@128572.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@128566.4]
  assign regs_121_clock = clock; // @[:@128575.4]
  assign regs_121_reset = io_reset; // @[:@128576.4 RegFile.scala 76:16:@128583.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@128582.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@128586.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@128580.4]
  assign regs_122_clock = clock; // @[:@128589.4]
  assign regs_122_reset = io_reset; // @[:@128590.4 RegFile.scala 76:16:@128597.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@128596.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@128600.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@128594.4]
  assign regs_123_clock = clock; // @[:@128603.4]
  assign regs_123_reset = io_reset; // @[:@128604.4 RegFile.scala 76:16:@128611.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@128610.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@128614.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@128608.4]
  assign regs_124_clock = clock; // @[:@128617.4]
  assign regs_124_reset = io_reset; // @[:@128618.4 RegFile.scala 76:16:@128625.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@128624.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@128628.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@128622.4]
  assign regs_125_clock = clock; // @[:@128631.4]
  assign regs_125_reset = io_reset; // @[:@128632.4 RegFile.scala 76:16:@128639.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@128638.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@128642.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@128636.4]
  assign regs_126_clock = clock; // @[:@128645.4]
  assign regs_126_reset = io_reset; // @[:@128646.4 RegFile.scala 76:16:@128653.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@128652.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@128656.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@128650.4]
  assign regs_127_clock = clock; // @[:@128659.4]
  assign regs_127_reset = io_reset; // @[:@128660.4 RegFile.scala 76:16:@128667.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@128666.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@128670.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@128664.4]
  assign regs_128_clock = clock; // @[:@128673.4]
  assign regs_128_reset = io_reset; // @[:@128674.4 RegFile.scala 76:16:@128681.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@128680.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@128684.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@128678.4]
  assign regs_129_clock = clock; // @[:@128687.4]
  assign regs_129_reset = io_reset; // @[:@128688.4 RegFile.scala 76:16:@128695.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@128694.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@128698.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@128692.4]
  assign regs_130_clock = clock; // @[:@128701.4]
  assign regs_130_reset = io_reset; // @[:@128702.4 RegFile.scala 76:16:@128709.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@128708.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@128712.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@128706.4]
  assign regs_131_clock = clock; // @[:@128715.4]
  assign regs_131_reset = io_reset; // @[:@128716.4 RegFile.scala 76:16:@128723.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@128722.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@128726.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@128720.4]
  assign regs_132_clock = clock; // @[:@128729.4]
  assign regs_132_reset = io_reset; // @[:@128730.4 RegFile.scala 76:16:@128737.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@128736.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@128740.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@128734.4]
  assign regs_133_clock = clock; // @[:@128743.4]
  assign regs_133_reset = io_reset; // @[:@128744.4 RegFile.scala 76:16:@128751.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@128750.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@128754.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@128748.4]
  assign regs_134_clock = clock; // @[:@128757.4]
  assign regs_134_reset = io_reset; // @[:@128758.4 RegFile.scala 76:16:@128765.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@128764.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@128768.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@128762.4]
  assign regs_135_clock = clock; // @[:@128771.4]
  assign regs_135_reset = io_reset; // @[:@128772.4 RegFile.scala 76:16:@128779.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@128778.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@128782.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@128776.4]
  assign regs_136_clock = clock; // @[:@128785.4]
  assign regs_136_reset = io_reset; // @[:@128786.4 RegFile.scala 76:16:@128793.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@128792.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@128796.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@128790.4]
  assign regs_137_clock = clock; // @[:@128799.4]
  assign regs_137_reset = io_reset; // @[:@128800.4 RegFile.scala 76:16:@128807.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@128806.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@128810.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@128804.4]
  assign regs_138_clock = clock; // @[:@128813.4]
  assign regs_138_reset = io_reset; // @[:@128814.4 RegFile.scala 76:16:@128821.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@128820.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@128824.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@128818.4]
  assign regs_139_clock = clock; // @[:@128827.4]
  assign regs_139_reset = io_reset; // @[:@128828.4 RegFile.scala 76:16:@128835.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@128834.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@128838.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@128832.4]
  assign regs_140_clock = clock; // @[:@128841.4]
  assign regs_140_reset = io_reset; // @[:@128842.4 RegFile.scala 76:16:@128849.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@128848.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@128852.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@128846.4]
  assign regs_141_clock = clock; // @[:@128855.4]
  assign regs_141_reset = io_reset; // @[:@128856.4 RegFile.scala 76:16:@128863.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@128862.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@128866.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@128860.4]
  assign regs_142_clock = clock; // @[:@128869.4]
  assign regs_142_reset = io_reset; // @[:@128870.4 RegFile.scala 76:16:@128877.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@128876.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@128880.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@128874.4]
  assign regs_143_clock = clock; // @[:@128883.4]
  assign regs_143_reset = io_reset; // @[:@128884.4 RegFile.scala 76:16:@128891.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@128890.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@128894.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@128888.4]
  assign regs_144_clock = clock; // @[:@128897.4]
  assign regs_144_reset = io_reset; // @[:@128898.4 RegFile.scala 76:16:@128905.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@128904.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@128908.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@128902.4]
  assign regs_145_clock = clock; // @[:@128911.4]
  assign regs_145_reset = io_reset; // @[:@128912.4 RegFile.scala 76:16:@128919.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@128918.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@128922.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@128916.4]
  assign regs_146_clock = clock; // @[:@128925.4]
  assign regs_146_reset = io_reset; // @[:@128926.4 RegFile.scala 76:16:@128933.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@128932.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@128936.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@128930.4]
  assign regs_147_clock = clock; // @[:@128939.4]
  assign regs_147_reset = io_reset; // @[:@128940.4 RegFile.scala 76:16:@128947.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@128946.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@128950.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@128944.4]
  assign regs_148_clock = clock; // @[:@128953.4]
  assign regs_148_reset = io_reset; // @[:@128954.4 RegFile.scala 76:16:@128961.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@128960.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@128964.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@128958.4]
  assign regs_149_clock = clock; // @[:@128967.4]
  assign regs_149_reset = io_reset; // @[:@128968.4 RegFile.scala 76:16:@128975.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@128974.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@128978.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@128972.4]
  assign regs_150_clock = clock; // @[:@128981.4]
  assign regs_150_reset = io_reset; // @[:@128982.4 RegFile.scala 76:16:@128989.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@128988.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@128992.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@128986.4]
  assign regs_151_clock = clock; // @[:@128995.4]
  assign regs_151_reset = io_reset; // @[:@128996.4 RegFile.scala 76:16:@129003.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@129002.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@129006.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@129000.4]
  assign regs_152_clock = clock; // @[:@129009.4]
  assign regs_152_reset = io_reset; // @[:@129010.4 RegFile.scala 76:16:@129017.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@129016.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@129020.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@129014.4]
  assign regs_153_clock = clock; // @[:@129023.4]
  assign regs_153_reset = io_reset; // @[:@129024.4 RegFile.scala 76:16:@129031.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@129030.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@129034.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@129028.4]
  assign regs_154_clock = clock; // @[:@129037.4]
  assign regs_154_reset = io_reset; // @[:@129038.4 RegFile.scala 76:16:@129045.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@129044.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@129048.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@129042.4]
  assign regs_155_clock = clock; // @[:@129051.4]
  assign regs_155_reset = io_reset; // @[:@129052.4 RegFile.scala 76:16:@129059.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@129058.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@129062.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@129056.4]
  assign regs_156_clock = clock; // @[:@129065.4]
  assign regs_156_reset = io_reset; // @[:@129066.4 RegFile.scala 76:16:@129073.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@129072.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@129076.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@129070.4]
  assign regs_157_clock = clock; // @[:@129079.4]
  assign regs_157_reset = io_reset; // @[:@129080.4 RegFile.scala 76:16:@129087.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@129086.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@129090.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@129084.4]
  assign regs_158_clock = clock; // @[:@129093.4]
  assign regs_158_reset = io_reset; // @[:@129094.4 RegFile.scala 76:16:@129101.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@129100.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@129104.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@129098.4]
  assign regs_159_clock = clock; // @[:@129107.4]
  assign regs_159_reset = io_reset; // @[:@129108.4 RegFile.scala 76:16:@129115.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@129114.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@129118.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@129112.4]
  assign regs_160_clock = clock; // @[:@129121.4]
  assign regs_160_reset = io_reset; // @[:@129122.4 RegFile.scala 76:16:@129129.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@129128.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@129132.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@129126.4]
  assign regs_161_clock = clock; // @[:@129135.4]
  assign regs_161_reset = io_reset; // @[:@129136.4 RegFile.scala 76:16:@129143.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@129142.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@129146.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@129140.4]
  assign regs_162_clock = clock; // @[:@129149.4]
  assign regs_162_reset = io_reset; // @[:@129150.4 RegFile.scala 76:16:@129157.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@129156.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@129160.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@129154.4]
  assign regs_163_clock = clock; // @[:@129163.4]
  assign regs_163_reset = io_reset; // @[:@129164.4 RegFile.scala 76:16:@129171.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@129170.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@129174.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@129168.4]
  assign regs_164_clock = clock; // @[:@129177.4]
  assign regs_164_reset = io_reset; // @[:@129178.4 RegFile.scala 76:16:@129185.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@129184.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@129188.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@129182.4]
  assign regs_165_clock = clock; // @[:@129191.4]
  assign regs_165_reset = io_reset; // @[:@129192.4 RegFile.scala 76:16:@129199.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@129198.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@129202.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@129196.4]
  assign regs_166_clock = clock; // @[:@129205.4]
  assign regs_166_reset = io_reset; // @[:@129206.4 RegFile.scala 76:16:@129213.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@129212.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@129216.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@129210.4]
  assign regs_167_clock = clock; // @[:@129219.4]
  assign regs_167_reset = io_reset; // @[:@129220.4 RegFile.scala 76:16:@129227.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@129226.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@129230.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@129224.4]
  assign regs_168_clock = clock; // @[:@129233.4]
  assign regs_168_reset = io_reset; // @[:@129234.4 RegFile.scala 76:16:@129241.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@129240.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@129244.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@129238.4]
  assign regs_169_clock = clock; // @[:@129247.4]
  assign regs_169_reset = io_reset; // @[:@129248.4 RegFile.scala 76:16:@129255.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@129254.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@129258.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@129252.4]
  assign regs_170_clock = clock; // @[:@129261.4]
  assign regs_170_reset = io_reset; // @[:@129262.4 RegFile.scala 76:16:@129269.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@129268.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@129272.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@129266.4]
  assign regs_171_clock = clock; // @[:@129275.4]
  assign regs_171_reset = io_reset; // @[:@129276.4 RegFile.scala 76:16:@129283.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@129282.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@129286.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@129280.4]
  assign regs_172_clock = clock; // @[:@129289.4]
  assign regs_172_reset = io_reset; // @[:@129290.4 RegFile.scala 76:16:@129297.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@129296.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@129300.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@129294.4]
  assign regs_173_clock = clock; // @[:@129303.4]
  assign regs_173_reset = io_reset; // @[:@129304.4 RegFile.scala 76:16:@129311.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@129310.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@129314.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@129308.4]
  assign regs_174_clock = clock; // @[:@129317.4]
  assign regs_174_reset = io_reset; // @[:@129318.4 RegFile.scala 76:16:@129325.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@129324.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@129328.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@129322.4]
  assign regs_175_clock = clock; // @[:@129331.4]
  assign regs_175_reset = io_reset; // @[:@129332.4 RegFile.scala 76:16:@129339.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@129338.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@129342.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@129336.4]
  assign regs_176_clock = clock; // @[:@129345.4]
  assign regs_176_reset = io_reset; // @[:@129346.4 RegFile.scala 76:16:@129353.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@129352.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@129356.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@129350.4]
  assign regs_177_clock = clock; // @[:@129359.4]
  assign regs_177_reset = io_reset; // @[:@129360.4 RegFile.scala 76:16:@129367.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@129366.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@129370.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@129364.4]
  assign regs_178_clock = clock; // @[:@129373.4]
  assign regs_178_reset = io_reset; // @[:@129374.4 RegFile.scala 76:16:@129381.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@129380.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@129384.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@129378.4]
  assign regs_179_clock = clock; // @[:@129387.4]
  assign regs_179_reset = io_reset; // @[:@129388.4 RegFile.scala 76:16:@129395.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@129394.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@129398.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@129392.4]
  assign regs_180_clock = clock; // @[:@129401.4]
  assign regs_180_reset = io_reset; // @[:@129402.4 RegFile.scala 76:16:@129409.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@129408.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@129412.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@129406.4]
  assign regs_181_clock = clock; // @[:@129415.4]
  assign regs_181_reset = io_reset; // @[:@129416.4 RegFile.scala 76:16:@129423.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@129422.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@129426.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@129420.4]
  assign regs_182_clock = clock; // @[:@129429.4]
  assign regs_182_reset = io_reset; // @[:@129430.4 RegFile.scala 76:16:@129437.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@129436.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@129440.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@129434.4]
  assign regs_183_clock = clock; // @[:@129443.4]
  assign regs_183_reset = io_reset; // @[:@129444.4 RegFile.scala 76:16:@129451.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@129450.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@129454.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@129448.4]
  assign regs_184_clock = clock; // @[:@129457.4]
  assign regs_184_reset = io_reset; // @[:@129458.4 RegFile.scala 76:16:@129465.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@129464.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@129468.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@129462.4]
  assign regs_185_clock = clock; // @[:@129471.4]
  assign regs_185_reset = io_reset; // @[:@129472.4 RegFile.scala 76:16:@129479.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@129478.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@129482.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@129476.4]
  assign regs_186_clock = clock; // @[:@129485.4]
  assign regs_186_reset = io_reset; // @[:@129486.4 RegFile.scala 76:16:@129493.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@129492.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@129496.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@129490.4]
  assign regs_187_clock = clock; // @[:@129499.4]
  assign regs_187_reset = io_reset; // @[:@129500.4 RegFile.scala 76:16:@129507.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@129506.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@129510.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@129504.4]
  assign regs_188_clock = clock; // @[:@129513.4]
  assign regs_188_reset = io_reset; // @[:@129514.4 RegFile.scala 76:16:@129521.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@129520.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@129524.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@129518.4]
  assign regs_189_clock = clock; // @[:@129527.4]
  assign regs_189_reset = io_reset; // @[:@129528.4 RegFile.scala 76:16:@129535.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@129534.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@129538.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@129532.4]
  assign regs_190_clock = clock; // @[:@129541.4]
  assign regs_190_reset = io_reset; // @[:@129542.4 RegFile.scala 76:16:@129549.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@129548.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@129552.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@129546.4]
  assign regs_191_clock = clock; // @[:@129555.4]
  assign regs_191_reset = io_reset; // @[:@129556.4 RegFile.scala 76:16:@129563.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@129562.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@129566.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@129560.4]
  assign regs_192_clock = clock; // @[:@129569.4]
  assign regs_192_reset = io_reset; // @[:@129570.4 RegFile.scala 76:16:@129577.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@129576.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@129580.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@129574.4]
  assign regs_193_clock = clock; // @[:@129583.4]
  assign regs_193_reset = io_reset; // @[:@129584.4 RegFile.scala 76:16:@129591.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@129590.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@129594.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@129588.4]
  assign regs_194_clock = clock; // @[:@129597.4]
  assign regs_194_reset = io_reset; // @[:@129598.4 RegFile.scala 76:16:@129605.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@129604.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@129608.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@129602.4]
  assign regs_195_clock = clock; // @[:@129611.4]
  assign regs_195_reset = io_reset; // @[:@129612.4 RegFile.scala 76:16:@129619.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@129618.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@129622.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@129616.4]
  assign regs_196_clock = clock; // @[:@129625.4]
  assign regs_196_reset = io_reset; // @[:@129626.4 RegFile.scala 76:16:@129633.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@129632.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@129636.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@129630.4]
  assign regs_197_clock = clock; // @[:@129639.4]
  assign regs_197_reset = io_reset; // @[:@129640.4 RegFile.scala 76:16:@129647.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@129646.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@129650.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@129644.4]
  assign regs_198_clock = clock; // @[:@129653.4]
  assign regs_198_reset = io_reset; // @[:@129654.4 RegFile.scala 76:16:@129661.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@129660.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@129664.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@129658.4]
  assign regs_199_clock = clock; // @[:@129667.4]
  assign regs_199_reset = io_reset; // @[:@129668.4 RegFile.scala 76:16:@129675.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@129674.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@129678.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@129672.4]
  assign regs_200_clock = clock; // @[:@129681.4]
  assign regs_200_reset = io_reset; // @[:@129682.4 RegFile.scala 76:16:@129689.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@129688.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@129692.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@129686.4]
  assign regs_201_clock = clock; // @[:@129695.4]
  assign regs_201_reset = io_reset; // @[:@129696.4 RegFile.scala 76:16:@129703.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@129702.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@129706.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@129700.4]
  assign regs_202_clock = clock; // @[:@129709.4]
  assign regs_202_reset = io_reset; // @[:@129710.4 RegFile.scala 76:16:@129717.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@129716.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@129720.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@129714.4]
  assign regs_203_clock = clock; // @[:@129723.4]
  assign regs_203_reset = io_reset; // @[:@129724.4 RegFile.scala 76:16:@129731.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@129730.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@129734.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@129728.4]
  assign regs_204_clock = clock; // @[:@129737.4]
  assign regs_204_reset = io_reset; // @[:@129738.4 RegFile.scala 76:16:@129745.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@129744.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@129748.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@129742.4]
  assign regs_205_clock = clock; // @[:@129751.4]
  assign regs_205_reset = io_reset; // @[:@129752.4 RegFile.scala 76:16:@129759.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@129758.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@129762.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@129756.4]
  assign regs_206_clock = clock; // @[:@129765.4]
  assign regs_206_reset = io_reset; // @[:@129766.4 RegFile.scala 76:16:@129773.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@129772.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@129776.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@129770.4]
  assign regs_207_clock = clock; // @[:@129779.4]
  assign regs_207_reset = io_reset; // @[:@129780.4 RegFile.scala 76:16:@129787.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@129786.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@129790.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@129784.4]
  assign regs_208_clock = clock; // @[:@129793.4]
  assign regs_208_reset = io_reset; // @[:@129794.4 RegFile.scala 76:16:@129801.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@129800.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@129804.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@129798.4]
  assign regs_209_clock = clock; // @[:@129807.4]
  assign regs_209_reset = io_reset; // @[:@129808.4 RegFile.scala 76:16:@129815.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@129814.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@129818.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@129812.4]
  assign regs_210_clock = clock; // @[:@129821.4]
  assign regs_210_reset = io_reset; // @[:@129822.4 RegFile.scala 76:16:@129829.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@129828.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@129832.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@129826.4]
  assign regs_211_clock = clock; // @[:@129835.4]
  assign regs_211_reset = io_reset; // @[:@129836.4 RegFile.scala 76:16:@129843.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@129842.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@129846.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@129840.4]
  assign regs_212_clock = clock; // @[:@129849.4]
  assign regs_212_reset = io_reset; // @[:@129850.4 RegFile.scala 76:16:@129857.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@129856.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@129860.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@129854.4]
  assign regs_213_clock = clock; // @[:@129863.4]
  assign regs_213_reset = io_reset; // @[:@129864.4 RegFile.scala 76:16:@129871.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@129870.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@129874.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@129868.4]
  assign regs_214_clock = clock; // @[:@129877.4]
  assign regs_214_reset = io_reset; // @[:@129878.4 RegFile.scala 76:16:@129885.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@129884.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@129888.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@129882.4]
  assign regs_215_clock = clock; // @[:@129891.4]
  assign regs_215_reset = io_reset; // @[:@129892.4 RegFile.scala 76:16:@129899.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@129898.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@129902.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@129896.4]
  assign regs_216_clock = clock; // @[:@129905.4]
  assign regs_216_reset = io_reset; // @[:@129906.4 RegFile.scala 76:16:@129913.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@129912.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@129916.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@129910.4]
  assign regs_217_clock = clock; // @[:@129919.4]
  assign regs_217_reset = io_reset; // @[:@129920.4 RegFile.scala 76:16:@129927.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@129926.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@129930.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@129924.4]
  assign regs_218_clock = clock; // @[:@129933.4]
  assign regs_218_reset = io_reset; // @[:@129934.4 RegFile.scala 76:16:@129941.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@129940.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@129944.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@129938.4]
  assign regs_219_clock = clock; // @[:@129947.4]
  assign regs_219_reset = io_reset; // @[:@129948.4 RegFile.scala 76:16:@129955.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@129954.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@129958.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@129952.4]
  assign regs_220_clock = clock; // @[:@129961.4]
  assign regs_220_reset = io_reset; // @[:@129962.4 RegFile.scala 76:16:@129969.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@129968.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@129972.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@129966.4]
  assign regs_221_clock = clock; // @[:@129975.4]
  assign regs_221_reset = io_reset; // @[:@129976.4 RegFile.scala 76:16:@129983.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@129982.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@129986.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@129980.4]
  assign regs_222_clock = clock; // @[:@129989.4]
  assign regs_222_reset = io_reset; // @[:@129990.4 RegFile.scala 76:16:@129997.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@129996.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@130000.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@129994.4]
  assign regs_223_clock = clock; // @[:@130003.4]
  assign regs_223_reset = io_reset; // @[:@130004.4 RegFile.scala 76:16:@130011.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@130010.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@130014.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@130008.4]
  assign regs_224_clock = clock; // @[:@130017.4]
  assign regs_224_reset = io_reset; // @[:@130018.4 RegFile.scala 76:16:@130025.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@130024.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@130028.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@130022.4]
  assign regs_225_clock = clock; // @[:@130031.4]
  assign regs_225_reset = io_reset; // @[:@130032.4 RegFile.scala 76:16:@130039.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@130038.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@130042.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@130036.4]
  assign regs_226_clock = clock; // @[:@130045.4]
  assign regs_226_reset = io_reset; // @[:@130046.4 RegFile.scala 76:16:@130053.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@130052.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@130056.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@130050.4]
  assign regs_227_clock = clock; // @[:@130059.4]
  assign regs_227_reset = io_reset; // @[:@130060.4 RegFile.scala 76:16:@130067.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@130066.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@130070.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@130064.4]
  assign regs_228_clock = clock; // @[:@130073.4]
  assign regs_228_reset = io_reset; // @[:@130074.4 RegFile.scala 76:16:@130081.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@130080.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@130084.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@130078.4]
  assign regs_229_clock = clock; // @[:@130087.4]
  assign regs_229_reset = io_reset; // @[:@130088.4 RegFile.scala 76:16:@130095.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@130094.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@130098.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@130092.4]
  assign regs_230_clock = clock; // @[:@130101.4]
  assign regs_230_reset = io_reset; // @[:@130102.4 RegFile.scala 76:16:@130109.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@130108.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@130112.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@130106.4]
  assign regs_231_clock = clock; // @[:@130115.4]
  assign regs_231_reset = io_reset; // @[:@130116.4 RegFile.scala 76:16:@130123.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@130122.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@130126.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@130120.4]
  assign regs_232_clock = clock; // @[:@130129.4]
  assign regs_232_reset = io_reset; // @[:@130130.4 RegFile.scala 76:16:@130137.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@130136.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@130140.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@130134.4]
  assign regs_233_clock = clock; // @[:@130143.4]
  assign regs_233_reset = io_reset; // @[:@130144.4 RegFile.scala 76:16:@130151.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@130150.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@130154.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@130148.4]
  assign regs_234_clock = clock; // @[:@130157.4]
  assign regs_234_reset = io_reset; // @[:@130158.4 RegFile.scala 76:16:@130165.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@130164.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@130168.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@130162.4]
  assign regs_235_clock = clock; // @[:@130171.4]
  assign regs_235_reset = io_reset; // @[:@130172.4 RegFile.scala 76:16:@130179.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@130178.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@130182.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@130176.4]
  assign regs_236_clock = clock; // @[:@130185.4]
  assign regs_236_reset = io_reset; // @[:@130186.4 RegFile.scala 76:16:@130193.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@130192.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@130196.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@130190.4]
  assign regs_237_clock = clock; // @[:@130199.4]
  assign regs_237_reset = io_reset; // @[:@130200.4 RegFile.scala 76:16:@130207.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@130206.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@130210.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@130204.4]
  assign regs_238_clock = clock; // @[:@130213.4]
  assign regs_238_reset = io_reset; // @[:@130214.4 RegFile.scala 76:16:@130221.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@130220.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@130224.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@130218.4]
  assign regs_239_clock = clock; // @[:@130227.4]
  assign regs_239_reset = io_reset; // @[:@130228.4 RegFile.scala 76:16:@130235.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@130234.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@130238.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@130232.4]
  assign regs_240_clock = clock; // @[:@130241.4]
  assign regs_240_reset = io_reset; // @[:@130242.4 RegFile.scala 76:16:@130249.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@130248.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@130252.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@130246.4]
  assign regs_241_clock = clock; // @[:@130255.4]
  assign regs_241_reset = io_reset; // @[:@130256.4 RegFile.scala 76:16:@130263.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@130262.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@130266.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@130260.4]
  assign regs_242_clock = clock; // @[:@130269.4]
  assign regs_242_reset = io_reset; // @[:@130270.4 RegFile.scala 76:16:@130277.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@130276.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@130280.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@130274.4]
  assign regs_243_clock = clock; // @[:@130283.4]
  assign regs_243_reset = io_reset; // @[:@130284.4 RegFile.scala 76:16:@130291.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@130290.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@130294.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@130288.4]
  assign regs_244_clock = clock; // @[:@130297.4]
  assign regs_244_reset = io_reset; // @[:@130298.4 RegFile.scala 76:16:@130305.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@130304.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@130308.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@130302.4]
  assign regs_245_clock = clock; // @[:@130311.4]
  assign regs_245_reset = io_reset; // @[:@130312.4 RegFile.scala 76:16:@130319.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@130318.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@130322.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@130316.4]
  assign regs_246_clock = clock; // @[:@130325.4]
  assign regs_246_reset = io_reset; // @[:@130326.4 RegFile.scala 76:16:@130333.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@130332.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@130336.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@130330.4]
  assign regs_247_clock = clock; // @[:@130339.4]
  assign regs_247_reset = io_reset; // @[:@130340.4 RegFile.scala 76:16:@130347.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@130346.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@130350.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@130344.4]
  assign regs_248_clock = clock; // @[:@130353.4]
  assign regs_248_reset = io_reset; // @[:@130354.4 RegFile.scala 76:16:@130361.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@130360.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@130364.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@130358.4]
  assign regs_249_clock = clock; // @[:@130367.4]
  assign regs_249_reset = io_reset; // @[:@130368.4 RegFile.scala 76:16:@130375.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@130374.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@130378.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@130372.4]
  assign regs_250_clock = clock; // @[:@130381.4]
  assign regs_250_reset = io_reset; // @[:@130382.4 RegFile.scala 76:16:@130389.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@130388.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@130392.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@130386.4]
  assign regs_251_clock = clock; // @[:@130395.4]
  assign regs_251_reset = io_reset; // @[:@130396.4 RegFile.scala 76:16:@130403.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@130402.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@130406.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@130400.4]
  assign regs_252_clock = clock; // @[:@130409.4]
  assign regs_252_reset = io_reset; // @[:@130410.4 RegFile.scala 76:16:@130417.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@130416.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@130420.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@130414.4]
  assign regs_253_clock = clock; // @[:@130423.4]
  assign regs_253_reset = io_reset; // @[:@130424.4 RegFile.scala 76:16:@130431.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@130430.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@130434.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@130428.4]
  assign regs_254_clock = clock; // @[:@130437.4]
  assign regs_254_reset = io_reset; // @[:@130438.4 RegFile.scala 76:16:@130445.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@130444.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@130448.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@130442.4]
  assign regs_255_clock = clock; // @[:@130451.4]
  assign regs_255_reset = io_reset; // @[:@130452.4 RegFile.scala 76:16:@130459.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@130458.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@130462.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@130456.4]
  assign regs_256_clock = clock; // @[:@130465.4]
  assign regs_256_reset = io_reset; // @[:@130466.4 RegFile.scala 76:16:@130473.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@130472.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@130476.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@130470.4]
  assign regs_257_clock = clock; // @[:@130479.4]
  assign regs_257_reset = io_reset; // @[:@130480.4 RegFile.scala 76:16:@130487.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@130486.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@130490.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@130484.4]
  assign regs_258_clock = clock; // @[:@130493.4]
  assign regs_258_reset = io_reset; // @[:@130494.4 RegFile.scala 76:16:@130501.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@130500.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@130504.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@130498.4]
  assign regs_259_clock = clock; // @[:@130507.4]
  assign regs_259_reset = io_reset; // @[:@130508.4 RegFile.scala 76:16:@130515.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@130514.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@130518.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@130512.4]
  assign regs_260_clock = clock; // @[:@130521.4]
  assign regs_260_reset = io_reset; // @[:@130522.4 RegFile.scala 76:16:@130529.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@130528.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@130532.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@130526.4]
  assign regs_261_clock = clock; // @[:@130535.4]
  assign regs_261_reset = io_reset; // @[:@130536.4 RegFile.scala 76:16:@130543.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@130542.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@130546.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@130540.4]
  assign regs_262_clock = clock; // @[:@130549.4]
  assign regs_262_reset = io_reset; // @[:@130550.4 RegFile.scala 76:16:@130557.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@130556.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@130560.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@130554.4]
  assign regs_263_clock = clock; // @[:@130563.4]
  assign regs_263_reset = io_reset; // @[:@130564.4 RegFile.scala 76:16:@130571.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@130570.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@130574.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@130568.4]
  assign regs_264_clock = clock; // @[:@130577.4]
  assign regs_264_reset = io_reset; // @[:@130578.4 RegFile.scala 76:16:@130585.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@130584.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@130588.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@130582.4]
  assign regs_265_clock = clock; // @[:@130591.4]
  assign regs_265_reset = io_reset; // @[:@130592.4 RegFile.scala 76:16:@130599.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@130598.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@130602.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@130596.4]
  assign regs_266_clock = clock; // @[:@130605.4]
  assign regs_266_reset = io_reset; // @[:@130606.4 RegFile.scala 76:16:@130613.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@130612.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@130616.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@130610.4]
  assign regs_267_clock = clock; // @[:@130619.4]
  assign regs_267_reset = io_reset; // @[:@130620.4 RegFile.scala 76:16:@130627.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@130626.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@130630.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@130624.4]
  assign regs_268_clock = clock; // @[:@130633.4]
  assign regs_268_reset = io_reset; // @[:@130634.4 RegFile.scala 76:16:@130641.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@130640.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@130644.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@130638.4]
  assign regs_269_clock = clock; // @[:@130647.4]
  assign regs_269_reset = io_reset; // @[:@130648.4 RegFile.scala 76:16:@130655.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@130654.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@130658.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@130652.4]
  assign regs_270_clock = clock; // @[:@130661.4]
  assign regs_270_reset = io_reset; // @[:@130662.4 RegFile.scala 76:16:@130669.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@130668.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@130672.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@130666.4]
  assign regs_271_clock = clock; // @[:@130675.4]
  assign regs_271_reset = io_reset; // @[:@130676.4 RegFile.scala 76:16:@130683.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@130682.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@130686.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@130680.4]
  assign regs_272_clock = clock; // @[:@130689.4]
  assign regs_272_reset = io_reset; // @[:@130690.4 RegFile.scala 76:16:@130697.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@130696.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@130700.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@130694.4]
  assign regs_273_clock = clock; // @[:@130703.4]
  assign regs_273_reset = io_reset; // @[:@130704.4 RegFile.scala 76:16:@130711.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@130710.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@130714.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@130708.4]
  assign regs_274_clock = clock; // @[:@130717.4]
  assign regs_274_reset = io_reset; // @[:@130718.4 RegFile.scala 76:16:@130725.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@130724.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@130728.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@130722.4]
  assign regs_275_clock = clock; // @[:@130731.4]
  assign regs_275_reset = io_reset; // @[:@130732.4 RegFile.scala 76:16:@130739.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@130738.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@130742.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@130736.4]
  assign regs_276_clock = clock; // @[:@130745.4]
  assign regs_276_reset = io_reset; // @[:@130746.4 RegFile.scala 76:16:@130753.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@130752.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@130756.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@130750.4]
  assign regs_277_clock = clock; // @[:@130759.4]
  assign regs_277_reset = io_reset; // @[:@130760.4 RegFile.scala 76:16:@130767.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@130766.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@130770.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@130764.4]
  assign regs_278_clock = clock; // @[:@130773.4]
  assign regs_278_reset = io_reset; // @[:@130774.4 RegFile.scala 76:16:@130781.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@130780.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@130784.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@130778.4]
  assign regs_279_clock = clock; // @[:@130787.4]
  assign regs_279_reset = io_reset; // @[:@130788.4 RegFile.scala 76:16:@130795.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@130794.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@130798.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@130792.4]
  assign regs_280_clock = clock; // @[:@130801.4]
  assign regs_280_reset = io_reset; // @[:@130802.4 RegFile.scala 76:16:@130809.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@130808.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@130812.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@130806.4]
  assign regs_281_clock = clock; // @[:@130815.4]
  assign regs_281_reset = io_reset; // @[:@130816.4 RegFile.scala 76:16:@130823.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@130822.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@130826.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@130820.4]
  assign regs_282_clock = clock; // @[:@130829.4]
  assign regs_282_reset = io_reset; // @[:@130830.4 RegFile.scala 76:16:@130837.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@130836.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@130840.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@130834.4]
  assign regs_283_clock = clock; // @[:@130843.4]
  assign regs_283_reset = io_reset; // @[:@130844.4 RegFile.scala 76:16:@130851.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@130850.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@130854.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@130848.4]
  assign regs_284_clock = clock; // @[:@130857.4]
  assign regs_284_reset = io_reset; // @[:@130858.4 RegFile.scala 76:16:@130865.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@130864.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@130868.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@130862.4]
  assign regs_285_clock = clock; // @[:@130871.4]
  assign regs_285_reset = io_reset; // @[:@130872.4 RegFile.scala 76:16:@130879.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@130878.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@130882.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@130876.4]
  assign regs_286_clock = clock; // @[:@130885.4]
  assign regs_286_reset = io_reset; // @[:@130886.4 RegFile.scala 76:16:@130893.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@130892.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@130896.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@130890.4]
  assign regs_287_clock = clock; // @[:@130899.4]
  assign regs_287_reset = io_reset; // @[:@130900.4 RegFile.scala 76:16:@130907.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@130906.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@130910.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@130904.4]
  assign regs_288_clock = clock; // @[:@130913.4]
  assign regs_288_reset = io_reset; // @[:@130914.4 RegFile.scala 76:16:@130921.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@130920.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@130924.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@130918.4]
  assign regs_289_clock = clock; // @[:@130927.4]
  assign regs_289_reset = io_reset; // @[:@130928.4 RegFile.scala 76:16:@130935.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@130934.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@130938.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@130932.4]
  assign regs_290_clock = clock; // @[:@130941.4]
  assign regs_290_reset = io_reset; // @[:@130942.4 RegFile.scala 76:16:@130949.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@130948.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@130952.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@130946.4]
  assign regs_291_clock = clock; // @[:@130955.4]
  assign regs_291_reset = io_reset; // @[:@130956.4 RegFile.scala 76:16:@130963.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@130962.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@130966.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@130960.4]
  assign regs_292_clock = clock; // @[:@130969.4]
  assign regs_292_reset = io_reset; // @[:@130970.4 RegFile.scala 76:16:@130977.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@130976.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@130980.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@130974.4]
  assign regs_293_clock = clock; // @[:@130983.4]
  assign regs_293_reset = io_reset; // @[:@130984.4 RegFile.scala 76:16:@130991.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@130990.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@130994.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@130988.4]
  assign regs_294_clock = clock; // @[:@130997.4]
  assign regs_294_reset = io_reset; // @[:@130998.4 RegFile.scala 76:16:@131005.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@131004.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@131008.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@131002.4]
  assign regs_295_clock = clock; // @[:@131011.4]
  assign regs_295_reset = io_reset; // @[:@131012.4 RegFile.scala 76:16:@131019.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@131018.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@131022.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@131016.4]
  assign regs_296_clock = clock; // @[:@131025.4]
  assign regs_296_reset = io_reset; // @[:@131026.4 RegFile.scala 76:16:@131033.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@131032.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@131036.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@131030.4]
  assign regs_297_clock = clock; // @[:@131039.4]
  assign regs_297_reset = io_reset; // @[:@131040.4 RegFile.scala 76:16:@131047.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@131046.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@131050.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@131044.4]
  assign regs_298_clock = clock; // @[:@131053.4]
  assign regs_298_reset = io_reset; // @[:@131054.4 RegFile.scala 76:16:@131061.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@131060.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@131064.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@131058.4]
  assign regs_299_clock = clock; // @[:@131067.4]
  assign regs_299_reset = io_reset; // @[:@131068.4 RegFile.scala 76:16:@131075.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@131074.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@131078.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@131072.4]
  assign regs_300_clock = clock; // @[:@131081.4]
  assign regs_300_reset = io_reset; // @[:@131082.4 RegFile.scala 76:16:@131089.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@131088.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@131092.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@131086.4]
  assign regs_301_clock = clock; // @[:@131095.4]
  assign regs_301_reset = io_reset; // @[:@131096.4 RegFile.scala 76:16:@131103.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@131102.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@131106.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@131100.4]
  assign regs_302_clock = clock; // @[:@131109.4]
  assign regs_302_reset = io_reset; // @[:@131110.4 RegFile.scala 76:16:@131117.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@131116.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@131120.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@131114.4]
  assign regs_303_clock = clock; // @[:@131123.4]
  assign regs_303_reset = io_reset; // @[:@131124.4 RegFile.scala 76:16:@131131.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@131130.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@131134.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@131128.4]
  assign regs_304_clock = clock; // @[:@131137.4]
  assign regs_304_reset = io_reset; // @[:@131138.4 RegFile.scala 76:16:@131145.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@131144.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@131148.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@131142.4]
  assign regs_305_clock = clock; // @[:@131151.4]
  assign regs_305_reset = io_reset; // @[:@131152.4 RegFile.scala 76:16:@131159.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@131158.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@131162.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@131156.4]
  assign regs_306_clock = clock; // @[:@131165.4]
  assign regs_306_reset = io_reset; // @[:@131166.4 RegFile.scala 76:16:@131173.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@131172.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@131176.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@131170.4]
  assign regs_307_clock = clock; // @[:@131179.4]
  assign regs_307_reset = io_reset; // @[:@131180.4 RegFile.scala 76:16:@131187.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@131186.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@131190.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@131184.4]
  assign regs_308_clock = clock; // @[:@131193.4]
  assign regs_308_reset = io_reset; // @[:@131194.4 RegFile.scala 76:16:@131201.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@131200.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@131204.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@131198.4]
  assign regs_309_clock = clock; // @[:@131207.4]
  assign regs_309_reset = io_reset; // @[:@131208.4 RegFile.scala 76:16:@131215.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@131214.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@131218.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@131212.4]
  assign regs_310_clock = clock; // @[:@131221.4]
  assign regs_310_reset = io_reset; // @[:@131222.4 RegFile.scala 76:16:@131229.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@131228.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@131232.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@131226.4]
  assign regs_311_clock = clock; // @[:@131235.4]
  assign regs_311_reset = io_reset; // @[:@131236.4 RegFile.scala 76:16:@131243.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@131242.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@131246.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@131240.4]
  assign regs_312_clock = clock; // @[:@131249.4]
  assign regs_312_reset = io_reset; // @[:@131250.4 RegFile.scala 76:16:@131257.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@131256.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@131260.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@131254.4]
  assign regs_313_clock = clock; // @[:@131263.4]
  assign regs_313_reset = io_reset; // @[:@131264.4 RegFile.scala 76:16:@131271.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@131270.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@131274.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@131268.4]
  assign regs_314_clock = clock; // @[:@131277.4]
  assign regs_314_reset = io_reset; // @[:@131278.4 RegFile.scala 76:16:@131285.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@131284.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@131288.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@131282.4]
  assign regs_315_clock = clock; // @[:@131291.4]
  assign regs_315_reset = io_reset; // @[:@131292.4 RegFile.scala 76:16:@131299.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@131298.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@131302.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@131296.4]
  assign regs_316_clock = clock; // @[:@131305.4]
  assign regs_316_reset = io_reset; // @[:@131306.4 RegFile.scala 76:16:@131313.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@131312.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@131316.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@131310.4]
  assign regs_317_clock = clock; // @[:@131319.4]
  assign regs_317_reset = io_reset; // @[:@131320.4 RegFile.scala 76:16:@131327.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@131326.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@131330.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@131324.4]
  assign regs_318_clock = clock; // @[:@131333.4]
  assign regs_318_reset = io_reset; // @[:@131334.4 RegFile.scala 76:16:@131341.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@131340.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@131344.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@131338.4]
  assign regs_319_clock = clock; // @[:@131347.4]
  assign regs_319_reset = io_reset; // @[:@131348.4 RegFile.scala 76:16:@131355.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@131354.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@131358.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@131352.4]
  assign regs_320_clock = clock; // @[:@131361.4]
  assign regs_320_reset = io_reset; // @[:@131362.4 RegFile.scala 76:16:@131369.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@131368.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@131372.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@131366.4]
  assign regs_321_clock = clock; // @[:@131375.4]
  assign regs_321_reset = io_reset; // @[:@131376.4 RegFile.scala 76:16:@131383.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@131382.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@131386.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@131380.4]
  assign regs_322_clock = clock; // @[:@131389.4]
  assign regs_322_reset = io_reset; // @[:@131390.4 RegFile.scala 76:16:@131397.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@131396.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@131400.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@131394.4]
  assign regs_323_clock = clock; // @[:@131403.4]
  assign regs_323_reset = io_reset; // @[:@131404.4 RegFile.scala 76:16:@131411.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@131410.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@131414.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@131408.4]
  assign regs_324_clock = clock; // @[:@131417.4]
  assign regs_324_reset = io_reset; // @[:@131418.4 RegFile.scala 76:16:@131425.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@131424.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@131428.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@131422.4]
  assign regs_325_clock = clock; // @[:@131431.4]
  assign regs_325_reset = io_reset; // @[:@131432.4 RegFile.scala 76:16:@131439.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@131438.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@131442.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@131436.4]
  assign regs_326_clock = clock; // @[:@131445.4]
  assign regs_326_reset = io_reset; // @[:@131446.4 RegFile.scala 76:16:@131453.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@131452.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@131456.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@131450.4]
  assign regs_327_clock = clock; // @[:@131459.4]
  assign regs_327_reset = io_reset; // @[:@131460.4 RegFile.scala 76:16:@131467.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@131466.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@131470.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@131464.4]
  assign regs_328_clock = clock; // @[:@131473.4]
  assign regs_328_reset = io_reset; // @[:@131474.4 RegFile.scala 76:16:@131481.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@131480.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@131484.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@131478.4]
  assign regs_329_clock = clock; // @[:@131487.4]
  assign regs_329_reset = io_reset; // @[:@131488.4 RegFile.scala 76:16:@131495.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@131494.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@131498.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@131492.4]
  assign regs_330_clock = clock; // @[:@131501.4]
  assign regs_330_reset = io_reset; // @[:@131502.4 RegFile.scala 76:16:@131509.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@131508.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@131512.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@131506.4]
  assign regs_331_clock = clock; // @[:@131515.4]
  assign regs_331_reset = io_reset; // @[:@131516.4 RegFile.scala 76:16:@131523.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@131522.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@131526.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@131520.4]
  assign regs_332_clock = clock; // @[:@131529.4]
  assign regs_332_reset = io_reset; // @[:@131530.4 RegFile.scala 76:16:@131537.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@131536.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@131540.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@131534.4]
  assign regs_333_clock = clock; // @[:@131543.4]
  assign regs_333_reset = io_reset; // @[:@131544.4 RegFile.scala 76:16:@131551.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@131550.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@131554.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@131548.4]
  assign regs_334_clock = clock; // @[:@131557.4]
  assign regs_334_reset = io_reset; // @[:@131558.4 RegFile.scala 76:16:@131565.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@131564.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@131568.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@131562.4]
  assign regs_335_clock = clock; // @[:@131571.4]
  assign regs_335_reset = io_reset; // @[:@131572.4 RegFile.scala 76:16:@131579.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@131578.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@131582.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@131576.4]
  assign regs_336_clock = clock; // @[:@131585.4]
  assign regs_336_reset = io_reset; // @[:@131586.4 RegFile.scala 76:16:@131593.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@131592.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@131596.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@131590.4]
  assign regs_337_clock = clock; // @[:@131599.4]
  assign regs_337_reset = io_reset; // @[:@131600.4 RegFile.scala 76:16:@131607.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@131606.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@131610.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@131604.4]
  assign regs_338_clock = clock; // @[:@131613.4]
  assign regs_338_reset = io_reset; // @[:@131614.4 RegFile.scala 76:16:@131621.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@131620.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@131624.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@131618.4]
  assign regs_339_clock = clock; // @[:@131627.4]
  assign regs_339_reset = io_reset; // @[:@131628.4 RegFile.scala 76:16:@131635.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@131634.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@131638.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@131632.4]
  assign regs_340_clock = clock; // @[:@131641.4]
  assign regs_340_reset = io_reset; // @[:@131642.4 RegFile.scala 76:16:@131649.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@131648.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@131652.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@131646.4]
  assign regs_341_clock = clock; // @[:@131655.4]
  assign regs_341_reset = io_reset; // @[:@131656.4 RegFile.scala 76:16:@131663.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@131662.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@131666.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@131660.4]
  assign regs_342_clock = clock; // @[:@131669.4]
  assign regs_342_reset = io_reset; // @[:@131670.4 RegFile.scala 76:16:@131677.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@131676.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@131680.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@131674.4]
  assign regs_343_clock = clock; // @[:@131683.4]
  assign regs_343_reset = io_reset; // @[:@131684.4 RegFile.scala 76:16:@131691.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@131690.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@131694.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@131688.4]
  assign regs_344_clock = clock; // @[:@131697.4]
  assign regs_344_reset = io_reset; // @[:@131698.4 RegFile.scala 76:16:@131705.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@131704.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@131708.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@131702.4]
  assign regs_345_clock = clock; // @[:@131711.4]
  assign regs_345_reset = io_reset; // @[:@131712.4 RegFile.scala 76:16:@131719.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@131718.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@131722.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@131716.4]
  assign regs_346_clock = clock; // @[:@131725.4]
  assign regs_346_reset = io_reset; // @[:@131726.4 RegFile.scala 76:16:@131733.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@131732.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@131736.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@131730.4]
  assign regs_347_clock = clock; // @[:@131739.4]
  assign regs_347_reset = io_reset; // @[:@131740.4 RegFile.scala 76:16:@131747.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@131746.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@131750.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@131744.4]
  assign regs_348_clock = clock; // @[:@131753.4]
  assign regs_348_reset = io_reset; // @[:@131754.4 RegFile.scala 76:16:@131761.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@131760.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@131764.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@131758.4]
  assign regs_349_clock = clock; // @[:@131767.4]
  assign regs_349_reset = io_reset; // @[:@131768.4 RegFile.scala 76:16:@131775.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@131774.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@131778.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@131772.4]
  assign regs_350_clock = clock; // @[:@131781.4]
  assign regs_350_reset = io_reset; // @[:@131782.4 RegFile.scala 76:16:@131789.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@131788.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@131792.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@131786.4]
  assign regs_351_clock = clock; // @[:@131795.4]
  assign regs_351_reset = io_reset; // @[:@131796.4 RegFile.scala 76:16:@131803.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@131802.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@131806.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@131800.4]
  assign regs_352_clock = clock; // @[:@131809.4]
  assign regs_352_reset = io_reset; // @[:@131810.4 RegFile.scala 76:16:@131817.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@131816.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@131820.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@131814.4]
  assign regs_353_clock = clock; // @[:@131823.4]
  assign regs_353_reset = io_reset; // @[:@131824.4 RegFile.scala 76:16:@131831.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@131830.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@131834.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@131828.4]
  assign regs_354_clock = clock; // @[:@131837.4]
  assign regs_354_reset = io_reset; // @[:@131838.4 RegFile.scala 76:16:@131845.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@131844.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@131848.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@131842.4]
  assign regs_355_clock = clock; // @[:@131851.4]
  assign regs_355_reset = io_reset; // @[:@131852.4 RegFile.scala 76:16:@131859.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@131858.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@131862.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@131856.4]
  assign regs_356_clock = clock; // @[:@131865.4]
  assign regs_356_reset = io_reset; // @[:@131866.4 RegFile.scala 76:16:@131873.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@131872.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@131876.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@131870.4]
  assign regs_357_clock = clock; // @[:@131879.4]
  assign regs_357_reset = io_reset; // @[:@131880.4 RegFile.scala 76:16:@131887.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@131886.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@131890.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@131884.4]
  assign regs_358_clock = clock; // @[:@131893.4]
  assign regs_358_reset = io_reset; // @[:@131894.4 RegFile.scala 76:16:@131901.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@131900.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@131904.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@131898.4]
  assign regs_359_clock = clock; // @[:@131907.4]
  assign regs_359_reset = io_reset; // @[:@131908.4 RegFile.scala 76:16:@131915.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@131914.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@131918.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@131912.4]
  assign regs_360_clock = clock; // @[:@131921.4]
  assign regs_360_reset = io_reset; // @[:@131922.4 RegFile.scala 76:16:@131929.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@131928.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@131932.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@131926.4]
  assign regs_361_clock = clock; // @[:@131935.4]
  assign regs_361_reset = io_reset; // @[:@131936.4 RegFile.scala 76:16:@131943.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@131942.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@131946.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@131940.4]
  assign regs_362_clock = clock; // @[:@131949.4]
  assign regs_362_reset = io_reset; // @[:@131950.4 RegFile.scala 76:16:@131957.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@131956.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@131960.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@131954.4]
  assign regs_363_clock = clock; // @[:@131963.4]
  assign regs_363_reset = io_reset; // @[:@131964.4 RegFile.scala 76:16:@131971.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@131970.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@131974.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@131968.4]
  assign regs_364_clock = clock; // @[:@131977.4]
  assign regs_364_reset = io_reset; // @[:@131978.4 RegFile.scala 76:16:@131985.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@131984.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@131988.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@131982.4]
  assign regs_365_clock = clock; // @[:@131991.4]
  assign regs_365_reset = io_reset; // @[:@131992.4 RegFile.scala 76:16:@131999.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@131998.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@132002.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@131996.4]
  assign regs_366_clock = clock; // @[:@132005.4]
  assign regs_366_reset = io_reset; // @[:@132006.4 RegFile.scala 76:16:@132013.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@132012.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@132016.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@132010.4]
  assign regs_367_clock = clock; // @[:@132019.4]
  assign regs_367_reset = io_reset; // @[:@132020.4 RegFile.scala 76:16:@132027.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@132026.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@132030.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@132024.4]
  assign regs_368_clock = clock; // @[:@132033.4]
  assign regs_368_reset = io_reset; // @[:@132034.4 RegFile.scala 76:16:@132041.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@132040.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@132044.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@132038.4]
  assign regs_369_clock = clock; // @[:@132047.4]
  assign regs_369_reset = io_reset; // @[:@132048.4 RegFile.scala 76:16:@132055.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@132054.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@132058.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@132052.4]
  assign regs_370_clock = clock; // @[:@132061.4]
  assign regs_370_reset = io_reset; // @[:@132062.4 RegFile.scala 76:16:@132069.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@132068.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@132072.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@132066.4]
  assign regs_371_clock = clock; // @[:@132075.4]
  assign regs_371_reset = io_reset; // @[:@132076.4 RegFile.scala 76:16:@132083.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@132082.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@132086.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@132080.4]
  assign regs_372_clock = clock; // @[:@132089.4]
  assign regs_372_reset = io_reset; // @[:@132090.4 RegFile.scala 76:16:@132097.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@132096.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@132100.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@132094.4]
  assign regs_373_clock = clock; // @[:@132103.4]
  assign regs_373_reset = io_reset; // @[:@132104.4 RegFile.scala 76:16:@132111.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@132110.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@132114.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@132108.4]
  assign regs_374_clock = clock; // @[:@132117.4]
  assign regs_374_reset = io_reset; // @[:@132118.4 RegFile.scala 76:16:@132125.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@132124.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@132128.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@132122.4]
  assign regs_375_clock = clock; // @[:@132131.4]
  assign regs_375_reset = io_reset; // @[:@132132.4 RegFile.scala 76:16:@132139.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@132138.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@132142.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@132136.4]
  assign regs_376_clock = clock; // @[:@132145.4]
  assign regs_376_reset = io_reset; // @[:@132146.4 RegFile.scala 76:16:@132153.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@132152.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@132156.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@132150.4]
  assign regs_377_clock = clock; // @[:@132159.4]
  assign regs_377_reset = io_reset; // @[:@132160.4 RegFile.scala 76:16:@132167.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@132166.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@132170.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@132164.4]
  assign regs_378_clock = clock; // @[:@132173.4]
  assign regs_378_reset = io_reset; // @[:@132174.4 RegFile.scala 76:16:@132181.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@132180.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@132184.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@132178.4]
  assign regs_379_clock = clock; // @[:@132187.4]
  assign regs_379_reset = io_reset; // @[:@132188.4 RegFile.scala 76:16:@132195.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@132194.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@132198.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@132192.4]
  assign regs_380_clock = clock; // @[:@132201.4]
  assign regs_380_reset = io_reset; // @[:@132202.4 RegFile.scala 76:16:@132209.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@132208.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@132212.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@132206.4]
  assign regs_381_clock = clock; // @[:@132215.4]
  assign regs_381_reset = io_reset; // @[:@132216.4 RegFile.scala 76:16:@132223.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@132222.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@132226.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@132220.4]
  assign regs_382_clock = clock; // @[:@132229.4]
  assign regs_382_reset = io_reset; // @[:@132230.4 RegFile.scala 76:16:@132237.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@132236.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@132240.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@132234.4]
  assign regs_383_clock = clock; // @[:@132243.4]
  assign regs_383_reset = io_reset; // @[:@132244.4 RegFile.scala 76:16:@132251.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@132250.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@132254.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@132248.4]
  assign regs_384_clock = clock; // @[:@132257.4]
  assign regs_384_reset = io_reset; // @[:@132258.4 RegFile.scala 76:16:@132265.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@132264.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@132268.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@132262.4]
  assign regs_385_clock = clock; // @[:@132271.4]
  assign regs_385_reset = io_reset; // @[:@132272.4 RegFile.scala 76:16:@132279.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@132278.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@132282.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@132276.4]
  assign regs_386_clock = clock; // @[:@132285.4]
  assign regs_386_reset = io_reset; // @[:@132286.4 RegFile.scala 76:16:@132293.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@132292.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@132296.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@132290.4]
  assign regs_387_clock = clock; // @[:@132299.4]
  assign regs_387_reset = io_reset; // @[:@132300.4 RegFile.scala 76:16:@132307.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@132306.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@132310.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@132304.4]
  assign regs_388_clock = clock; // @[:@132313.4]
  assign regs_388_reset = io_reset; // @[:@132314.4 RegFile.scala 76:16:@132321.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@132320.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@132324.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@132318.4]
  assign regs_389_clock = clock; // @[:@132327.4]
  assign regs_389_reset = io_reset; // @[:@132328.4 RegFile.scala 76:16:@132335.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@132334.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@132338.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@132332.4]
  assign regs_390_clock = clock; // @[:@132341.4]
  assign regs_390_reset = io_reset; // @[:@132342.4 RegFile.scala 76:16:@132349.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@132348.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@132352.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@132346.4]
  assign regs_391_clock = clock; // @[:@132355.4]
  assign regs_391_reset = io_reset; // @[:@132356.4 RegFile.scala 76:16:@132363.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@132362.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@132366.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@132360.4]
  assign regs_392_clock = clock; // @[:@132369.4]
  assign regs_392_reset = io_reset; // @[:@132370.4 RegFile.scala 76:16:@132377.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@132376.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@132380.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@132374.4]
  assign regs_393_clock = clock; // @[:@132383.4]
  assign regs_393_reset = io_reset; // @[:@132384.4 RegFile.scala 76:16:@132391.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@132390.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@132394.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@132388.4]
  assign regs_394_clock = clock; // @[:@132397.4]
  assign regs_394_reset = io_reset; // @[:@132398.4 RegFile.scala 76:16:@132405.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@132404.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@132408.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@132402.4]
  assign regs_395_clock = clock; // @[:@132411.4]
  assign regs_395_reset = io_reset; // @[:@132412.4 RegFile.scala 76:16:@132419.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@132418.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@132422.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@132416.4]
  assign regs_396_clock = clock; // @[:@132425.4]
  assign regs_396_reset = io_reset; // @[:@132426.4 RegFile.scala 76:16:@132433.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@132432.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@132436.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@132430.4]
  assign regs_397_clock = clock; // @[:@132439.4]
  assign regs_397_reset = io_reset; // @[:@132440.4 RegFile.scala 76:16:@132447.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@132446.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@132450.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@132444.4]
  assign regs_398_clock = clock; // @[:@132453.4]
  assign regs_398_reset = io_reset; // @[:@132454.4 RegFile.scala 76:16:@132461.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@132460.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@132464.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@132458.4]
  assign regs_399_clock = clock; // @[:@132467.4]
  assign regs_399_reset = io_reset; // @[:@132468.4 RegFile.scala 76:16:@132475.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@132474.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@132478.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@132472.4]
  assign regs_400_clock = clock; // @[:@132481.4]
  assign regs_400_reset = io_reset; // @[:@132482.4 RegFile.scala 76:16:@132489.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@132488.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@132492.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@132486.4]
  assign regs_401_clock = clock; // @[:@132495.4]
  assign regs_401_reset = io_reset; // @[:@132496.4 RegFile.scala 76:16:@132503.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@132502.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@132506.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@132500.4]
  assign regs_402_clock = clock; // @[:@132509.4]
  assign regs_402_reset = io_reset; // @[:@132510.4 RegFile.scala 76:16:@132517.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@132516.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@132520.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@132514.4]
  assign regs_403_clock = clock; // @[:@132523.4]
  assign regs_403_reset = io_reset; // @[:@132524.4 RegFile.scala 76:16:@132531.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@132530.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@132534.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@132528.4]
  assign regs_404_clock = clock; // @[:@132537.4]
  assign regs_404_reset = io_reset; // @[:@132538.4 RegFile.scala 76:16:@132545.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@132544.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@132548.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@132542.4]
  assign regs_405_clock = clock; // @[:@132551.4]
  assign regs_405_reset = io_reset; // @[:@132552.4 RegFile.scala 76:16:@132559.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@132558.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@132562.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@132556.4]
  assign regs_406_clock = clock; // @[:@132565.4]
  assign regs_406_reset = io_reset; // @[:@132566.4 RegFile.scala 76:16:@132573.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@132572.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@132576.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@132570.4]
  assign regs_407_clock = clock; // @[:@132579.4]
  assign regs_407_reset = io_reset; // @[:@132580.4 RegFile.scala 76:16:@132587.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@132586.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@132590.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@132584.4]
  assign regs_408_clock = clock; // @[:@132593.4]
  assign regs_408_reset = io_reset; // @[:@132594.4 RegFile.scala 76:16:@132601.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@132600.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@132604.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@132598.4]
  assign regs_409_clock = clock; // @[:@132607.4]
  assign regs_409_reset = io_reset; // @[:@132608.4 RegFile.scala 76:16:@132615.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@132614.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@132618.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@132612.4]
  assign regs_410_clock = clock; // @[:@132621.4]
  assign regs_410_reset = io_reset; // @[:@132622.4 RegFile.scala 76:16:@132629.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@132628.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@132632.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@132626.4]
  assign regs_411_clock = clock; // @[:@132635.4]
  assign regs_411_reset = io_reset; // @[:@132636.4 RegFile.scala 76:16:@132643.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@132642.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@132646.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@132640.4]
  assign regs_412_clock = clock; // @[:@132649.4]
  assign regs_412_reset = io_reset; // @[:@132650.4 RegFile.scala 76:16:@132657.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@132656.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@132660.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@132654.4]
  assign regs_413_clock = clock; // @[:@132663.4]
  assign regs_413_reset = io_reset; // @[:@132664.4 RegFile.scala 76:16:@132671.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@132670.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@132674.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@132668.4]
  assign regs_414_clock = clock; // @[:@132677.4]
  assign regs_414_reset = io_reset; // @[:@132678.4 RegFile.scala 76:16:@132685.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@132684.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@132688.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@132682.4]
  assign regs_415_clock = clock; // @[:@132691.4]
  assign regs_415_reset = io_reset; // @[:@132692.4 RegFile.scala 76:16:@132699.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@132698.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@132702.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@132696.4]
  assign regs_416_clock = clock; // @[:@132705.4]
  assign regs_416_reset = io_reset; // @[:@132706.4 RegFile.scala 76:16:@132713.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@132712.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@132716.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@132710.4]
  assign regs_417_clock = clock; // @[:@132719.4]
  assign regs_417_reset = io_reset; // @[:@132720.4 RegFile.scala 76:16:@132727.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@132726.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@132730.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@132724.4]
  assign regs_418_clock = clock; // @[:@132733.4]
  assign regs_418_reset = io_reset; // @[:@132734.4 RegFile.scala 76:16:@132741.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@132740.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@132744.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@132738.4]
  assign regs_419_clock = clock; // @[:@132747.4]
  assign regs_419_reset = io_reset; // @[:@132748.4 RegFile.scala 76:16:@132755.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@132754.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@132758.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@132752.4]
  assign regs_420_clock = clock; // @[:@132761.4]
  assign regs_420_reset = io_reset; // @[:@132762.4 RegFile.scala 76:16:@132769.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@132768.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@132772.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@132766.4]
  assign regs_421_clock = clock; // @[:@132775.4]
  assign regs_421_reset = io_reset; // @[:@132776.4 RegFile.scala 76:16:@132783.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@132782.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@132786.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@132780.4]
  assign regs_422_clock = clock; // @[:@132789.4]
  assign regs_422_reset = io_reset; // @[:@132790.4 RegFile.scala 76:16:@132797.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@132796.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@132800.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@132794.4]
  assign regs_423_clock = clock; // @[:@132803.4]
  assign regs_423_reset = io_reset; // @[:@132804.4 RegFile.scala 76:16:@132811.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@132810.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@132814.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@132808.4]
  assign regs_424_clock = clock; // @[:@132817.4]
  assign regs_424_reset = io_reset; // @[:@132818.4 RegFile.scala 76:16:@132825.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@132824.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@132828.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@132822.4]
  assign regs_425_clock = clock; // @[:@132831.4]
  assign regs_425_reset = io_reset; // @[:@132832.4 RegFile.scala 76:16:@132839.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@132838.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@132842.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@132836.4]
  assign regs_426_clock = clock; // @[:@132845.4]
  assign regs_426_reset = io_reset; // @[:@132846.4 RegFile.scala 76:16:@132853.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@132852.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@132856.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@132850.4]
  assign regs_427_clock = clock; // @[:@132859.4]
  assign regs_427_reset = io_reset; // @[:@132860.4 RegFile.scala 76:16:@132867.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@132866.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@132870.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@132864.4]
  assign regs_428_clock = clock; // @[:@132873.4]
  assign regs_428_reset = io_reset; // @[:@132874.4 RegFile.scala 76:16:@132881.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@132880.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@132884.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@132878.4]
  assign regs_429_clock = clock; // @[:@132887.4]
  assign regs_429_reset = io_reset; // @[:@132888.4 RegFile.scala 76:16:@132895.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@132894.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@132898.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@132892.4]
  assign regs_430_clock = clock; // @[:@132901.4]
  assign regs_430_reset = io_reset; // @[:@132902.4 RegFile.scala 76:16:@132909.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@132908.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@132912.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@132906.4]
  assign regs_431_clock = clock; // @[:@132915.4]
  assign regs_431_reset = io_reset; // @[:@132916.4 RegFile.scala 76:16:@132923.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@132922.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@132926.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@132920.4]
  assign regs_432_clock = clock; // @[:@132929.4]
  assign regs_432_reset = io_reset; // @[:@132930.4 RegFile.scala 76:16:@132937.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@132936.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@132940.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@132934.4]
  assign regs_433_clock = clock; // @[:@132943.4]
  assign regs_433_reset = io_reset; // @[:@132944.4 RegFile.scala 76:16:@132951.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@132950.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@132954.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@132948.4]
  assign regs_434_clock = clock; // @[:@132957.4]
  assign regs_434_reset = io_reset; // @[:@132958.4 RegFile.scala 76:16:@132965.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@132964.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@132968.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@132962.4]
  assign regs_435_clock = clock; // @[:@132971.4]
  assign regs_435_reset = io_reset; // @[:@132972.4 RegFile.scala 76:16:@132979.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@132978.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@132982.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@132976.4]
  assign regs_436_clock = clock; // @[:@132985.4]
  assign regs_436_reset = io_reset; // @[:@132986.4 RegFile.scala 76:16:@132993.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@132992.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@132996.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@132990.4]
  assign regs_437_clock = clock; // @[:@132999.4]
  assign regs_437_reset = io_reset; // @[:@133000.4 RegFile.scala 76:16:@133007.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@133006.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@133010.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@133004.4]
  assign regs_438_clock = clock; // @[:@133013.4]
  assign regs_438_reset = io_reset; // @[:@133014.4 RegFile.scala 76:16:@133021.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@133020.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@133024.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@133018.4]
  assign regs_439_clock = clock; // @[:@133027.4]
  assign regs_439_reset = io_reset; // @[:@133028.4 RegFile.scala 76:16:@133035.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@133034.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@133038.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@133032.4]
  assign regs_440_clock = clock; // @[:@133041.4]
  assign regs_440_reset = io_reset; // @[:@133042.4 RegFile.scala 76:16:@133049.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@133048.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@133052.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@133046.4]
  assign regs_441_clock = clock; // @[:@133055.4]
  assign regs_441_reset = io_reset; // @[:@133056.4 RegFile.scala 76:16:@133063.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@133062.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@133066.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@133060.4]
  assign regs_442_clock = clock; // @[:@133069.4]
  assign regs_442_reset = io_reset; // @[:@133070.4 RegFile.scala 76:16:@133077.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@133076.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@133080.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@133074.4]
  assign regs_443_clock = clock; // @[:@133083.4]
  assign regs_443_reset = io_reset; // @[:@133084.4 RegFile.scala 76:16:@133091.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@133090.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@133094.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@133088.4]
  assign regs_444_clock = clock; // @[:@133097.4]
  assign regs_444_reset = io_reset; // @[:@133098.4 RegFile.scala 76:16:@133105.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@133104.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@133108.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@133102.4]
  assign regs_445_clock = clock; // @[:@133111.4]
  assign regs_445_reset = io_reset; // @[:@133112.4 RegFile.scala 76:16:@133119.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@133118.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@133122.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@133116.4]
  assign regs_446_clock = clock; // @[:@133125.4]
  assign regs_446_reset = io_reset; // @[:@133126.4 RegFile.scala 76:16:@133133.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@133132.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@133136.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@133130.4]
  assign regs_447_clock = clock; // @[:@133139.4]
  assign regs_447_reset = io_reset; // @[:@133140.4 RegFile.scala 76:16:@133147.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@133146.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@133150.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@133144.4]
  assign regs_448_clock = clock; // @[:@133153.4]
  assign regs_448_reset = io_reset; // @[:@133154.4 RegFile.scala 76:16:@133161.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@133160.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@133164.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@133158.4]
  assign regs_449_clock = clock; // @[:@133167.4]
  assign regs_449_reset = io_reset; // @[:@133168.4 RegFile.scala 76:16:@133175.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@133174.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@133178.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@133172.4]
  assign regs_450_clock = clock; // @[:@133181.4]
  assign regs_450_reset = io_reset; // @[:@133182.4 RegFile.scala 76:16:@133189.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@133188.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@133192.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@133186.4]
  assign regs_451_clock = clock; // @[:@133195.4]
  assign regs_451_reset = io_reset; // @[:@133196.4 RegFile.scala 76:16:@133203.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@133202.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@133206.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@133200.4]
  assign regs_452_clock = clock; // @[:@133209.4]
  assign regs_452_reset = io_reset; // @[:@133210.4 RegFile.scala 76:16:@133217.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@133216.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@133220.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@133214.4]
  assign regs_453_clock = clock; // @[:@133223.4]
  assign regs_453_reset = io_reset; // @[:@133224.4 RegFile.scala 76:16:@133231.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@133230.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@133234.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@133228.4]
  assign regs_454_clock = clock; // @[:@133237.4]
  assign regs_454_reset = io_reset; // @[:@133238.4 RegFile.scala 76:16:@133245.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@133244.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@133248.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@133242.4]
  assign regs_455_clock = clock; // @[:@133251.4]
  assign regs_455_reset = io_reset; // @[:@133252.4 RegFile.scala 76:16:@133259.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@133258.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@133262.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@133256.4]
  assign regs_456_clock = clock; // @[:@133265.4]
  assign regs_456_reset = io_reset; // @[:@133266.4 RegFile.scala 76:16:@133273.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@133272.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@133276.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@133270.4]
  assign regs_457_clock = clock; // @[:@133279.4]
  assign regs_457_reset = io_reset; // @[:@133280.4 RegFile.scala 76:16:@133287.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@133286.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@133290.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@133284.4]
  assign regs_458_clock = clock; // @[:@133293.4]
  assign regs_458_reset = io_reset; // @[:@133294.4 RegFile.scala 76:16:@133301.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@133300.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@133304.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@133298.4]
  assign regs_459_clock = clock; // @[:@133307.4]
  assign regs_459_reset = io_reset; // @[:@133308.4 RegFile.scala 76:16:@133315.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@133314.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@133318.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@133312.4]
  assign regs_460_clock = clock; // @[:@133321.4]
  assign regs_460_reset = io_reset; // @[:@133322.4 RegFile.scala 76:16:@133329.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@133328.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@133332.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@133326.4]
  assign regs_461_clock = clock; // @[:@133335.4]
  assign regs_461_reset = io_reset; // @[:@133336.4 RegFile.scala 76:16:@133343.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@133342.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@133346.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@133340.4]
  assign regs_462_clock = clock; // @[:@133349.4]
  assign regs_462_reset = io_reset; // @[:@133350.4 RegFile.scala 76:16:@133357.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@133356.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@133360.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@133354.4]
  assign regs_463_clock = clock; // @[:@133363.4]
  assign regs_463_reset = io_reset; // @[:@133364.4 RegFile.scala 76:16:@133371.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@133370.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@133374.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@133368.4]
  assign regs_464_clock = clock; // @[:@133377.4]
  assign regs_464_reset = io_reset; // @[:@133378.4 RegFile.scala 76:16:@133385.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@133384.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@133388.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@133382.4]
  assign regs_465_clock = clock; // @[:@133391.4]
  assign regs_465_reset = io_reset; // @[:@133392.4 RegFile.scala 76:16:@133399.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@133398.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@133402.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@133396.4]
  assign regs_466_clock = clock; // @[:@133405.4]
  assign regs_466_reset = io_reset; // @[:@133406.4 RegFile.scala 76:16:@133413.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@133412.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@133416.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@133410.4]
  assign regs_467_clock = clock; // @[:@133419.4]
  assign regs_467_reset = io_reset; // @[:@133420.4 RegFile.scala 76:16:@133427.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@133426.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@133430.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@133424.4]
  assign regs_468_clock = clock; // @[:@133433.4]
  assign regs_468_reset = io_reset; // @[:@133434.4 RegFile.scala 76:16:@133441.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@133440.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@133444.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@133438.4]
  assign regs_469_clock = clock; // @[:@133447.4]
  assign regs_469_reset = io_reset; // @[:@133448.4 RegFile.scala 76:16:@133455.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@133454.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@133458.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@133452.4]
  assign regs_470_clock = clock; // @[:@133461.4]
  assign regs_470_reset = io_reset; // @[:@133462.4 RegFile.scala 76:16:@133469.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@133468.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@133472.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@133466.4]
  assign regs_471_clock = clock; // @[:@133475.4]
  assign regs_471_reset = io_reset; // @[:@133476.4 RegFile.scala 76:16:@133483.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@133482.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@133486.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@133480.4]
  assign regs_472_clock = clock; // @[:@133489.4]
  assign regs_472_reset = io_reset; // @[:@133490.4 RegFile.scala 76:16:@133497.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@133496.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@133500.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@133494.4]
  assign regs_473_clock = clock; // @[:@133503.4]
  assign regs_473_reset = io_reset; // @[:@133504.4 RegFile.scala 76:16:@133511.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@133510.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@133514.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@133508.4]
  assign regs_474_clock = clock; // @[:@133517.4]
  assign regs_474_reset = io_reset; // @[:@133518.4 RegFile.scala 76:16:@133525.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@133524.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@133528.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@133522.4]
  assign regs_475_clock = clock; // @[:@133531.4]
  assign regs_475_reset = io_reset; // @[:@133532.4 RegFile.scala 76:16:@133539.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@133538.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@133542.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@133536.4]
  assign regs_476_clock = clock; // @[:@133545.4]
  assign regs_476_reset = io_reset; // @[:@133546.4 RegFile.scala 76:16:@133553.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@133552.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@133556.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@133550.4]
  assign regs_477_clock = clock; // @[:@133559.4]
  assign regs_477_reset = io_reset; // @[:@133560.4 RegFile.scala 76:16:@133567.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@133566.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@133570.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@133564.4]
  assign regs_478_clock = clock; // @[:@133573.4]
  assign regs_478_reset = io_reset; // @[:@133574.4 RegFile.scala 76:16:@133581.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@133580.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@133584.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@133578.4]
  assign regs_479_clock = clock; // @[:@133587.4]
  assign regs_479_reset = io_reset; // @[:@133588.4 RegFile.scala 76:16:@133595.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@133594.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@133598.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@133592.4]
  assign regs_480_clock = clock; // @[:@133601.4]
  assign regs_480_reset = io_reset; // @[:@133602.4 RegFile.scala 76:16:@133609.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@133608.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@133612.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@133606.4]
  assign regs_481_clock = clock; // @[:@133615.4]
  assign regs_481_reset = io_reset; // @[:@133616.4 RegFile.scala 76:16:@133623.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@133622.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@133626.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@133620.4]
  assign regs_482_clock = clock; // @[:@133629.4]
  assign regs_482_reset = io_reset; // @[:@133630.4 RegFile.scala 76:16:@133637.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@133636.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@133640.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@133634.4]
  assign regs_483_clock = clock; // @[:@133643.4]
  assign regs_483_reset = io_reset; // @[:@133644.4 RegFile.scala 76:16:@133651.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@133650.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@133654.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@133648.4]
  assign regs_484_clock = clock; // @[:@133657.4]
  assign regs_484_reset = io_reset; // @[:@133658.4 RegFile.scala 76:16:@133665.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@133664.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@133668.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@133662.4]
  assign regs_485_clock = clock; // @[:@133671.4]
  assign regs_485_reset = io_reset; // @[:@133672.4 RegFile.scala 76:16:@133679.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@133678.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@133682.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@133676.4]
  assign regs_486_clock = clock; // @[:@133685.4]
  assign regs_486_reset = io_reset; // @[:@133686.4 RegFile.scala 76:16:@133693.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@133692.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@133696.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@133690.4]
  assign regs_487_clock = clock; // @[:@133699.4]
  assign regs_487_reset = io_reset; // @[:@133700.4 RegFile.scala 76:16:@133707.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@133706.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@133710.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@133704.4]
  assign regs_488_clock = clock; // @[:@133713.4]
  assign regs_488_reset = io_reset; // @[:@133714.4 RegFile.scala 76:16:@133721.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@133720.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@133724.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@133718.4]
  assign regs_489_clock = clock; // @[:@133727.4]
  assign regs_489_reset = io_reset; // @[:@133728.4 RegFile.scala 76:16:@133735.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@133734.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@133738.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@133732.4]
  assign regs_490_clock = clock; // @[:@133741.4]
  assign regs_490_reset = io_reset; // @[:@133742.4 RegFile.scala 76:16:@133749.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@133748.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@133752.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@133746.4]
  assign regs_491_clock = clock; // @[:@133755.4]
  assign regs_491_reset = io_reset; // @[:@133756.4 RegFile.scala 76:16:@133763.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@133762.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@133766.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@133760.4]
  assign regs_492_clock = clock; // @[:@133769.4]
  assign regs_492_reset = io_reset; // @[:@133770.4 RegFile.scala 76:16:@133777.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@133776.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@133780.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@133774.4]
  assign regs_493_clock = clock; // @[:@133783.4]
  assign regs_493_reset = io_reset; // @[:@133784.4 RegFile.scala 76:16:@133791.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@133790.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@133794.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@133788.4]
  assign regs_494_clock = clock; // @[:@133797.4]
  assign regs_494_reset = io_reset; // @[:@133798.4 RegFile.scala 76:16:@133805.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@133804.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@133808.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@133802.4]
  assign regs_495_clock = clock; // @[:@133811.4]
  assign regs_495_reset = io_reset; // @[:@133812.4 RegFile.scala 76:16:@133819.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@133818.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@133822.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@133816.4]
  assign regs_496_clock = clock; // @[:@133825.4]
  assign regs_496_reset = io_reset; // @[:@133826.4 RegFile.scala 76:16:@133833.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@133832.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@133836.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@133830.4]
  assign regs_497_clock = clock; // @[:@133839.4]
  assign regs_497_reset = io_reset; // @[:@133840.4 RegFile.scala 76:16:@133847.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@133846.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@133850.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@133844.4]
  assign regs_498_clock = clock; // @[:@133853.4]
  assign regs_498_reset = io_reset; // @[:@133854.4 RegFile.scala 76:16:@133861.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@133860.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@133864.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@133858.4]
  assign regs_499_clock = clock; // @[:@133867.4]
  assign regs_499_reset = io_reset; // @[:@133868.4 RegFile.scala 76:16:@133875.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@133874.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@133878.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@133872.4]
  assign regs_500_clock = clock; // @[:@133881.4]
  assign regs_500_reset = io_reset; // @[:@133882.4 RegFile.scala 76:16:@133889.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@133888.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@133892.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@133886.4]
  assign regs_501_clock = clock; // @[:@133895.4]
  assign regs_501_reset = io_reset; // @[:@133896.4 RegFile.scala 76:16:@133903.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@133902.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@133906.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@133900.4]
  assign regs_502_clock = clock; // @[:@133909.4]
  assign regs_502_reset = io_reset; // @[:@133910.4 RegFile.scala 76:16:@133917.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@133916.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@133920.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@133914.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@134429.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@134430.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@134431.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@134432.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@134433.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@134434.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@134435.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@134436.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@134437.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@134438.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@134439.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@134440.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@134441.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@134442.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@134443.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@134444.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@134445.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@134446.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@134447.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@134448.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@134449.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@134450.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@134451.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@134452.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@134453.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@134454.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@134455.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@134456.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@134457.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@134458.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@134459.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@134460.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@134461.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@134462.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@134463.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@134464.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@134465.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@134466.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@134467.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@134468.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@134469.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@134470.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@134471.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@134472.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@134473.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@134474.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@134475.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@134476.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@134477.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@134478.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@134479.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@134480.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@134481.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@134482.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@134483.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@134484.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@134485.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@134486.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@134487.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@134488.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@134489.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@134490.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@134491.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@134492.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@134493.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@134494.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@134495.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@134496.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@134497.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@134498.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@134499.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@134500.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@134501.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@134502.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@134503.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@134504.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@134505.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@134506.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@134507.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@134508.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@134509.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@134510.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@134511.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@134512.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@134513.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@134514.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@134515.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@134516.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@134517.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@134518.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@134519.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@134520.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@134521.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@134522.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@134523.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@134524.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@134525.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@134526.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@134527.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@134528.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@134529.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@134530.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@134531.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@134532.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@134533.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@134534.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@134535.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@134536.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@134537.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@134538.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@134539.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@134540.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@134541.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@134542.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@134543.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@134544.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@134545.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@134546.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@134547.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@134548.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@134549.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@134550.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@134551.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@134552.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@134553.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@134554.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@134555.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@134556.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@134557.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@134558.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@134559.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@134560.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@134561.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@134562.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@134563.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@134564.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@134565.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@134566.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@134567.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@134568.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@134569.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@134570.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@134571.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@134572.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@134573.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@134574.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@134575.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@134576.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@134577.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@134578.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@134579.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@134580.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@134581.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@134582.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@134583.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@134584.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@134585.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@134586.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@134587.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@134588.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@134589.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@134590.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@134591.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@134592.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@134593.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@134594.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@134595.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@134596.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@134597.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@134598.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@134599.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@134600.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@134601.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@134602.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@134603.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@134604.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@134605.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@134606.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@134607.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@134608.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@134609.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@134610.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@134611.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@134612.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@134613.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@134614.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@134615.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@134616.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@134617.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@134618.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@134619.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@134620.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@134621.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@134622.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@134623.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@134624.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@134625.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@134626.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@134627.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@134628.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@134629.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@134630.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@134631.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@134632.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@134633.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@134634.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@134635.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@134636.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@134637.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@134638.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@134639.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@134640.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@134641.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@134642.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@134643.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@134644.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@134645.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@134646.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@134647.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@134648.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@134649.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@134650.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@134651.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@134652.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@134653.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@134654.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@134655.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@134656.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@134657.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@134658.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@134659.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@134660.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@134661.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@134662.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@134663.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@134664.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@134665.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@134666.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@134667.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@134668.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@134669.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@134670.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@134671.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@134672.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@134673.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@134674.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@134675.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@134676.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@134677.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@134678.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@134679.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@134680.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@134681.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@134682.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@134683.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@134684.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@134685.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@134686.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@134687.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@134688.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@134689.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@134690.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@134691.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@134692.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@134693.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@134694.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@134695.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@134696.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@134697.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@134698.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@134699.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@134700.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@134701.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@134702.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@134703.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@134704.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@134705.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@134706.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@134707.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@134708.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@134709.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@134710.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@134711.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@134712.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@134713.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@134714.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@134715.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@134716.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@134717.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@134718.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@134719.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@134720.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@134721.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@134722.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@134723.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@134724.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@134725.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@134726.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@134727.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@134728.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@134729.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@134730.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@134731.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@134732.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@134733.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@134734.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@134735.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@134736.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@134737.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@134738.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@134739.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@134740.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@134741.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@134742.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@134743.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@134744.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@134745.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@134746.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@134747.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@134748.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@134749.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@134750.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@134751.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@134752.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@134753.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@134754.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@134755.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@134756.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@134757.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@134758.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@134759.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@134760.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@134761.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@134762.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@134763.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@134764.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@134765.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@134766.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@134767.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@134768.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@134769.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@134770.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@134771.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@134772.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@134773.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@134774.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@134775.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@134776.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@134777.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@134778.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@134779.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@134780.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@134781.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@134782.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@134783.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@134784.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@134785.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@134786.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@134787.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@134788.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@134789.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@134790.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@134791.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@134792.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@134793.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@134794.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@134795.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@134796.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@134797.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@134798.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@134799.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@134800.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@134801.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@134802.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@134803.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@134804.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@134805.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@134806.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@134807.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@134808.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@134809.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@134810.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@134811.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@134812.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@134813.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@134814.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@134815.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@134816.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@134817.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@134818.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@134819.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@134820.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@134821.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@134822.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@134823.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@134824.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@134825.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@134826.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@134827.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@134828.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@134829.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@134830.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@134831.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@134832.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@134833.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@134834.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@134835.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@134836.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@134837.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@134838.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@134839.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@134840.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@134841.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@134842.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@134843.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@134844.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@134845.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@134846.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@134847.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@134848.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@134849.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@134850.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@134851.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@134852.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@134853.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@134854.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@134855.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@134856.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@134857.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@134858.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@134859.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@134860.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@134861.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@134862.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@134863.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@134864.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@134865.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@134866.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@134867.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@134868.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@134869.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@134870.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@134871.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@134872.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@134873.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@134874.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@134875.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@134876.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@134877.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@134878.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@134879.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@134880.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@134881.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@134882.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@134883.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@134884.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@134885.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@134886.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@134887.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@134888.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@134889.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@134890.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@134891.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@134892.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@134893.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@134894.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@134895.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@134896.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@134897.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@134898.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@134899.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@134900.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@134901.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@134902.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@134903.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@134904.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@134905.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@134906.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@134907.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@134908.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@134909.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@134910.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@134911.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@134912.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@134913.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@134914.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@134915.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@134916.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@134917.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@134918.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@134919.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@134920.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@134921.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@134922.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@134923.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@134924.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@134925.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@134926.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@134927.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@134928.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@134929.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@134930.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@134931.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@134932.4]
endmodule
module RetimeWrapper_826( // @[:@134956.2]
  input         clock, // @[:@134957.4]
  input         reset, // @[:@134958.4]
  input  [39:0] io_in, // @[:@134959.4]
  output [39:0] io_out // @[:@134959.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@134961.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@134961.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@134961.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@134961.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@134961.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@134961.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@134961.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@134974.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@134973.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@134972.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@134971.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@134970.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@134968.4]
endmodule
module FringeFF_503( // @[:@134976.2]
  input         clock, // @[:@134977.4]
  input         reset, // @[:@134978.4]
  input  [39:0] io_in, // @[:@134979.4]
  output [39:0] io_out, // @[:@134979.4]
  input         io_enable // @[:@134979.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@134982.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@134982.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@134982.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@134982.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@134987.4 package.scala 96:25:@134988.4]
  RetimeWrapper_826 RetimeWrapper ( // @[package.scala 93:22:@134982.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@134987.4 package.scala 96:25:@134988.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@134999.4]
  assign RetimeWrapper_clock = clock; // @[:@134983.4]
  assign RetimeWrapper_reset = reset; // @[:@134984.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@134985.4]
endmodule
module FringeCounter( // @[:@135001.2]
  input   clock, // @[:@135002.4]
  input   reset, // @[:@135003.4]
  input   io_enable, // @[:@135004.4]
  output  io_done // @[:@135004.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@135006.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@135006.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@135006.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@135006.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@135006.4]
  wire [40:0] count; // @[Cat.scala 30:58:@135013.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@135014.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@135015.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@135016.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@135018.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@135006.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@135013.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@135014.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@135015.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@135016.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@135018.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@135029.4]
  assign reg$_clock = clock; // @[:@135007.4]
  assign reg$_reset = reset; // @[:@135008.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@135020.6 FringeCounter.scala 37:15:@135023.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@135011.4]
endmodule
module FringeFF_504( // @[:@135063.2]
  input   clock, // @[:@135064.4]
  input   reset, // @[:@135065.4]
  input   io_in, // @[:@135066.4]
  input   io_reset, // @[:@135066.4]
  output  io_out, // @[:@135066.4]
  input   io_enable // @[:@135066.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@135069.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@135069.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@135069.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@135069.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@135069.4]
  wire  _T_18; // @[package.scala 96:25:@135074.4 package.scala 96:25:@135075.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@135080.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@135069.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@135074.4 package.scala 96:25:@135075.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@135080.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@135086.4]
  assign RetimeWrapper_clock = clock; // @[:@135070.4]
  assign RetimeWrapper_reset = reset; // @[:@135071.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@135073.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@135072.4]
endmodule
module Depulser( // @[:@135088.2]
  input   clock, // @[:@135089.4]
  input   reset, // @[:@135090.4]
  input   io_in, // @[:@135091.4]
  input   io_rst, // @[:@135091.4]
  output  io_out // @[:@135091.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@135093.4]
  wire  r_reset; // @[Depulser.scala 14:17:@135093.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@135093.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@135093.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@135093.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@135093.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@135093.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@135102.4]
  assign r_clock = clock; // @[:@135094.4]
  assign r_reset = reset; // @[:@135095.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@135097.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@135101.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@135100.4]
endmodule
module Fringe( // @[:@135104.2]
  input         clock, // @[:@135105.4]
  input         reset, // @[:@135106.4]
  input  [31:0] io_raddr, // @[:@135107.4]
  input         io_wen, // @[:@135107.4]
  input  [31:0] io_waddr, // @[:@135107.4]
  input  [63:0] io_wdata, // @[:@135107.4]
  output [63:0] io_rdata, // @[:@135107.4]
  output        io_enable, // @[:@135107.4]
  input         io_done, // @[:@135107.4]
  output        io_reset, // @[:@135107.4]
  output [63:0] io_argIns_0, // @[:@135107.4]
  output [63:0] io_argIns_1, // @[:@135107.4]
  input         io_argOuts_0_valid, // @[:@135107.4]
  input  [63:0] io_argOuts_0_bits, // @[:@135107.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@135107.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@135107.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@135107.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@135107.4]
  output        io_memStreams_stores_0_data_ready, // @[:@135107.4]
  input         io_memStreams_stores_0_data_valid, // @[:@135107.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@135107.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@135107.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@135107.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@135107.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@135107.4]
  input         io_dram_0_cmd_ready, // @[:@135107.4]
  output        io_dram_0_cmd_valid, // @[:@135107.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@135107.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@135107.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@135107.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@135107.4]
  input         io_dram_0_wdata_ready, // @[:@135107.4]
  output        io_dram_0_wdata_valid, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@135107.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@135107.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@135107.4]
  output        io_dram_0_rresp_ready, // @[:@135107.4]
  output        io_dram_0_wresp_ready, // @[:@135107.4]
  input         io_dram_0_wresp_valid, // @[:@135107.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@135107.4]
  input         io_dram_1_cmd_ready, // @[:@135107.4]
  output        io_dram_1_cmd_valid, // @[:@135107.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@135107.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@135107.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@135107.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@135107.4]
  input         io_dram_1_wdata_ready, // @[:@135107.4]
  output        io_dram_1_wdata_valid, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@135107.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@135107.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@135107.4]
  output        io_dram_1_rresp_ready, // @[:@135107.4]
  output        io_dram_1_wresp_ready, // @[:@135107.4]
  input         io_dram_1_wresp_valid, // @[:@135107.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@135107.4]
  input         io_dram_2_cmd_ready, // @[:@135107.4]
  output        io_dram_2_cmd_valid, // @[:@135107.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@135107.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@135107.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@135107.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@135107.4]
  input         io_dram_2_wdata_ready, // @[:@135107.4]
  output        io_dram_2_wdata_valid, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@135107.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@135107.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@135107.4]
  output        io_dram_2_rresp_ready, // @[:@135107.4]
  output        io_dram_2_wresp_ready, // @[:@135107.4]
  input         io_dram_2_wresp_valid, // @[:@135107.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@135107.4]
  input         io_dram_3_cmd_ready, // @[:@135107.4]
  output        io_dram_3_cmd_valid, // @[:@135107.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@135107.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@135107.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@135107.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@135107.4]
  input         io_dram_3_wdata_ready, // @[:@135107.4]
  output        io_dram_3_wdata_valid, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@135107.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@135107.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@135107.4]
  output        io_dram_3_rresp_ready, // @[:@135107.4]
  output        io_dram_3_wresp_ready, // @[:@135107.4]
  input         io_dram_3_wresp_valid, // @[:@135107.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@135107.4]
  input         io_heap_0_req_valid, // @[:@135107.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@135107.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@135107.4]
  output        io_heap_0_resp_valid, // @[:@135107.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@135107.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@135107.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@135113.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@135113.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@135113.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@135113.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@136106.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@136106.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@136106.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@137066.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@137066.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@137066.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@138026.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@138026.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@138026.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@138026.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@138986.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@138986.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@138986.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@138986.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@138986.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@138986.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@138986.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@138986.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@138986.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@138986.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@138986.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@138986.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@138995.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@138995.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@138995.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@138995.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@138995.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@138995.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@138995.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@138995.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@138995.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@141045.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@141045.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@141045.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@141045.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@141064.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@141064.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@141064.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@141064.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@141064.4]
  wire [63:0] _T_1020; // @[:@141022.4 :@141023.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@141024.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@141026.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@141028.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@141030.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@141032.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@141034.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@141036.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@141072.4]
  reg  _T_1047; // @[package.scala 152:20:@141075.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@141077.4]
  wire  _T_1049; // @[package.scala 153:8:@141078.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@141082.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@141083.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@141086.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@141087.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@141089.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@141090.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@141092.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@141095.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@141074.4 Fringe.scala 163:24:@141093.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@141074.4 Fringe.scala 162:28:@141091.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@141096.4]
  wire  alloc; // @[Fringe.scala 202:38:@142726.4]
  wire  dealloc; // @[Fringe.scala 203:40:@142727.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@142728.4]
  reg  _T_1572; // @[package.scala 152:20:@142729.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@142731.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@135113.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@136106.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@137066.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@138026.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@138986.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@138995.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@141045.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@141064.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@141022.4 :@141023.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@141024.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@141026.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@141028.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@141030.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@141032.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@141034.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@141036.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@141072.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@141077.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@141078.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@141082.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@141083.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@141086.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@141087.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@141089.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@141090.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@141092.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@141095.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@141074.4 Fringe.scala 163:24:@141093.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@141074.4 Fringe.scala 162:28:@141091.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@141096.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@142726.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@142727.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@142728.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@142731.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@141020.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@141040.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@141041.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@141062.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@141063.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@136032.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@136028.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@136023.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@136022.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142224.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142223.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142222.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142220.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142219.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142217.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142201.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142202.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142203.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142204.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142205.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142206.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142207.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142208.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142209.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142210.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142211.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142212.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142213.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142214.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142215.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142216.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142137.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142138.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142139.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142140.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142141.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142142.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142143.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142144.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142145.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142146.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142147.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142148.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142149.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142150.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142151.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142152.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142153.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142154.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142155.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142156.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142157.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142158.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142159.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142160.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142161.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142162.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142163.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142164.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142165.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142166.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142167.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142168.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142169.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142170.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142171.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142172.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142173.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142174.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142175.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142176.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142177.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142178.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142179.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142180.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142181.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142182.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142183.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142184.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142185.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142186.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142187.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142188.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142189.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142190.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142191.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142192.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142193.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142194.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142195.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142196.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142197.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142198.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142199.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142200.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142136.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142135.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142116.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142336.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142335.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142334.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142332.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142331.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142329.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142313.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142314.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142315.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142316.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142317.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142318.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142319.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142320.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142321.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142322.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142323.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142324.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142325.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142326.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142327.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142328.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142249.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142250.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142251.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142252.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142253.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142254.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142255.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142256.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142257.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142258.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142259.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142260.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142261.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142262.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142263.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142264.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142265.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142266.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142267.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142268.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142269.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142270.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142271.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142272.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142273.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142274.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142275.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142276.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142277.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142278.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142279.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142280.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142281.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142282.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142283.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142284.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142285.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142286.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142287.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142288.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142289.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142290.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142291.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142292.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142293.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142294.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142295.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142296.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142297.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142298.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142299.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142300.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142301.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142302.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142303.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142304.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142305.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142306.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142307.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142308.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142309.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142310.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142311.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142312.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142248.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142247.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142228.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142448.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142447.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142446.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142444.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142443.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142441.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142425.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142426.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142427.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142428.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142429.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142430.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142431.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142432.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142433.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142434.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142435.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142436.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142437.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142438.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142439.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142440.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142361.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142362.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142363.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142364.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142365.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142366.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142367.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142368.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142369.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142370.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142371.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142372.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142373.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142374.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142375.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142376.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142377.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142378.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142379.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142380.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142381.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142382.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142383.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142384.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142385.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142386.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142387.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142388.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142389.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142390.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142391.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142392.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142393.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142394.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142395.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142396.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142397.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142398.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142399.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142400.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142401.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142402.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142403.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142404.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142405.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142406.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142407.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142408.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142409.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142410.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142411.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142412.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142413.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142414.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142415.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142416.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142417.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142418.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142419.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142420.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142421.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142422.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142423.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142424.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142360.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142359.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142340.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142560.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142559.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142558.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142556.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142555.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142553.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142537.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142538.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142539.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142540.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142541.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142542.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142543.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142544.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142545.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142546.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142547.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142548.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142549.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142550.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142551.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142552.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142473.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142474.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142475.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142476.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142477.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142478.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142479.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142480.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142481.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142482.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142483.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142484.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142485.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142486.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142487.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142488.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142489.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142490.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142491.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142492.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142493.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142494.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142495.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142496.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142497.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142498.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142499.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142500.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142501.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142502.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142503.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142504.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142505.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142506.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142507.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142508.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142509.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142510.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142511.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142512.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142513.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142514.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142515.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142516.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142517.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142518.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142519.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142520.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142521.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142522.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142523.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142524.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142525.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142526.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142527.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142528.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142529.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142530.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142531.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142532.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142533.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142534.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142535.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142536.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142472.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142471.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142452.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@138991.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@138990.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@138989.4]
  assign dramArbs_0_clock = clock; // @[:@135114.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@135115.4 Fringe.scala 187:30:@142106.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142110.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@136031.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@136030.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@136029.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@136027.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@136026.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@136025.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@136024.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@142225.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@142218.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@142115.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@142114.4]
  assign dramArbs_1_clock = clock; // @[:@136107.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@136108.4 Fringe.scala 187:30:@142107.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142111.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@142337.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@142330.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@142227.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@142226.4]
  assign dramArbs_2_clock = clock; // @[:@137067.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@137068.4 Fringe.scala 187:30:@142108.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142112.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@142449.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@142442.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@142339.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@142338.4]
  assign dramArbs_3_clock = clock; // @[:@138027.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@138028.4 Fringe.scala 187:30:@142109.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142113.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@142561.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@142554.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@142451.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@142450.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@138994.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@138993.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@138992.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@142733.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@142734.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@142735.4]
  assign regs_clock = clock; // @[:@138996.4]
  assign regs_reset = reset; // @[:@138997.4 Fringe.scala 139:14:@141044.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@141016.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@141018.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@141017.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@141019.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@141042.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@141094.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@141098.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@141101.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@141100.4]
  assign timeoutCtr_clock = clock; // @[:@141046.4]
  assign timeoutCtr_reset = reset; // @[:@141047.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@141061.4]
  assign depulser_clock = clock; // @[:@141065.4]
  assign depulser_reset = reset; // @[:@141066.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@141071.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@141073.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@142750.2]
  input         clock, // @[:@142751.4]
  input         reset, // @[:@142752.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@142753.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@142753.4]
  input         io_S_AXI_AWVALID, // @[:@142753.4]
  output        io_S_AXI_AWREADY, // @[:@142753.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@142753.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@142753.4]
  input         io_S_AXI_ARVALID, // @[:@142753.4]
  output        io_S_AXI_ARREADY, // @[:@142753.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@142753.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@142753.4]
  input         io_S_AXI_WVALID, // @[:@142753.4]
  output        io_S_AXI_WREADY, // @[:@142753.4]
  output [31:0] io_S_AXI_RDATA, // @[:@142753.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@142753.4]
  output        io_S_AXI_RVALID, // @[:@142753.4]
  input         io_S_AXI_RREADY, // @[:@142753.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@142753.4]
  output        io_S_AXI_BVALID, // @[:@142753.4]
  input         io_S_AXI_BREADY, // @[:@142753.4]
  output [31:0] io_raddr, // @[:@142753.4]
  output        io_wen, // @[:@142753.4]
  output [31:0] io_waddr, // @[:@142753.4]
  output [31:0] io_wdata, // @[:@142753.4]
  input  [31:0] io_rdata // @[:@142753.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@142755.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142779.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142775.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142771.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@142770.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@142769.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142768.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@142766.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142765.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@142787.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@142790.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@142788.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@142789.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@142791.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@142786.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@142783.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@142782.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@142781.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142780.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@142778.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@142777.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142776.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@142774.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@142773.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142772.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142767.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142764.4]
endmodule
module MAGToAXI4Bridge( // @[:@142793.2]
  output         io_in_cmd_ready, // @[:@142796.4]
  input          io_in_cmd_valid, // @[:@142796.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@142796.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@142796.4]
  input          io_in_cmd_bits_isWr, // @[:@142796.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@142796.4]
  output         io_in_wdata_ready, // @[:@142796.4]
  input          io_in_wdata_valid, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@142796.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@142796.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@142796.4]
  input          io_in_wdata_bits_wlast, // @[:@142796.4]
  input          io_in_rresp_ready, // @[:@142796.4]
  input          io_in_wresp_ready, // @[:@142796.4]
  output         io_in_wresp_valid, // @[:@142796.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@142796.4]
  output [31:0]  io_M_AXI_AWID, // @[:@142796.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@142796.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@142796.4]
  output         io_M_AXI_AWVALID, // @[:@142796.4]
  input          io_M_AXI_AWREADY, // @[:@142796.4]
  output [31:0]  io_M_AXI_ARID, // @[:@142796.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@142796.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@142796.4]
  output         io_M_AXI_ARVALID, // @[:@142796.4]
  input          io_M_AXI_ARREADY, // @[:@142796.4]
  output [511:0] io_M_AXI_WDATA, // @[:@142796.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@142796.4]
  output         io_M_AXI_WLAST, // @[:@142796.4]
  output         io_M_AXI_WVALID, // @[:@142796.4]
  input          io_M_AXI_WREADY, // @[:@142796.4]
  output         io_M_AXI_RREADY, // @[:@142796.4]
  input  [31:0]  io_M_AXI_BID, // @[:@142796.4]
  input          io_M_AXI_BVALID, // @[:@142796.4]
  output         io_M_AXI_BREADY // @[:@142796.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@142953.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@142954.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@142955.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@142963.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@142990.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@142995.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@143006.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@143015.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@143024.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@143033.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@143042.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@143051.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@143059.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@142953.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@142954.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@142955.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@142963.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@142990.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@142995.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@143006.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@143015.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@143024.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@143033.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@143042.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@143051.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@143059.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@142967.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@143064.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@143117.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@143119.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@142968.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@142969.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@142973.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@142981.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@142951.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@142952.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@142956.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@142965.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@142997.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@143061.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@143062.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@143063.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@143114.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@143115.4]
endmodule
module FringeZynq( // @[:@144105.2]
  input          clock, // @[:@144106.4]
  input          reset, // @[:@144107.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@144108.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@144108.4]
  input          io_S_AXI_AWVALID, // @[:@144108.4]
  output         io_S_AXI_AWREADY, // @[:@144108.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@144108.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@144108.4]
  input          io_S_AXI_ARVALID, // @[:@144108.4]
  output         io_S_AXI_ARREADY, // @[:@144108.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@144108.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@144108.4]
  input          io_S_AXI_WVALID, // @[:@144108.4]
  output         io_S_AXI_WREADY, // @[:@144108.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@144108.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@144108.4]
  output         io_S_AXI_RVALID, // @[:@144108.4]
  input          io_S_AXI_RREADY, // @[:@144108.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@144108.4]
  output         io_S_AXI_BVALID, // @[:@144108.4]
  input          io_S_AXI_BREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@144108.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@144108.4]
  output         io_M_AXI_0_AWVALID, // @[:@144108.4]
  input          io_M_AXI_0_AWREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@144108.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@144108.4]
  output         io_M_AXI_0_ARVALID, // @[:@144108.4]
  input          io_M_AXI_0_ARREADY, // @[:@144108.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@144108.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@144108.4]
  output         io_M_AXI_0_WLAST, // @[:@144108.4]
  output         io_M_AXI_0_WVALID, // @[:@144108.4]
  input          io_M_AXI_0_WREADY, // @[:@144108.4]
  output         io_M_AXI_0_RREADY, // @[:@144108.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@144108.4]
  input          io_M_AXI_0_BVALID, // @[:@144108.4]
  output         io_M_AXI_0_BREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@144108.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@144108.4]
  output         io_M_AXI_1_AWVALID, // @[:@144108.4]
  input          io_M_AXI_1_AWREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@144108.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@144108.4]
  output         io_M_AXI_1_ARVALID, // @[:@144108.4]
  input          io_M_AXI_1_ARREADY, // @[:@144108.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@144108.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@144108.4]
  output         io_M_AXI_1_WLAST, // @[:@144108.4]
  output         io_M_AXI_1_WVALID, // @[:@144108.4]
  input          io_M_AXI_1_WREADY, // @[:@144108.4]
  output         io_M_AXI_1_RREADY, // @[:@144108.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@144108.4]
  input          io_M_AXI_1_BVALID, // @[:@144108.4]
  output         io_M_AXI_1_BREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@144108.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@144108.4]
  output         io_M_AXI_2_AWVALID, // @[:@144108.4]
  input          io_M_AXI_2_AWREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@144108.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@144108.4]
  output         io_M_AXI_2_ARVALID, // @[:@144108.4]
  input          io_M_AXI_2_ARREADY, // @[:@144108.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@144108.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@144108.4]
  output         io_M_AXI_2_WLAST, // @[:@144108.4]
  output         io_M_AXI_2_WVALID, // @[:@144108.4]
  input          io_M_AXI_2_WREADY, // @[:@144108.4]
  output         io_M_AXI_2_RREADY, // @[:@144108.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@144108.4]
  input          io_M_AXI_2_BVALID, // @[:@144108.4]
  output         io_M_AXI_2_BREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@144108.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@144108.4]
  output         io_M_AXI_3_AWVALID, // @[:@144108.4]
  input          io_M_AXI_3_AWREADY, // @[:@144108.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@144108.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@144108.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@144108.4]
  output         io_M_AXI_3_ARVALID, // @[:@144108.4]
  input          io_M_AXI_3_ARREADY, // @[:@144108.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@144108.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@144108.4]
  output         io_M_AXI_3_WLAST, // @[:@144108.4]
  output         io_M_AXI_3_WVALID, // @[:@144108.4]
  input          io_M_AXI_3_WREADY, // @[:@144108.4]
  output         io_M_AXI_3_RREADY, // @[:@144108.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@144108.4]
  input          io_M_AXI_3_BVALID, // @[:@144108.4]
  output         io_M_AXI_3_BREADY, // @[:@144108.4]
  output         io_enable, // @[:@144108.4]
  input          io_done, // @[:@144108.4]
  output         io_reset, // @[:@144108.4]
  output [63:0]  io_argIns_0, // @[:@144108.4]
  output [63:0]  io_argIns_1, // @[:@144108.4]
  input          io_argOuts_0_valid, // @[:@144108.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@144108.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@144108.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@144108.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@144108.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@144108.4]
  output         io_memStreams_stores_0_data_ready, // @[:@144108.4]
  input          io_memStreams_stores_0_data_valid, // @[:@144108.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@144108.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@144108.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@144108.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@144108.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@144108.4]
  input          io_heap_0_req_valid, // @[:@144108.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@144108.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@144108.4]
  output         io_heap_0_resp_valid, // @[:@144108.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@144108.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@144108.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@144579.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@144579.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@144579.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@145485.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@145485.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@145485.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@145485.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@145485.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@145485.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@145485.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@145485.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@145635.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@145635.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@145635.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@145635.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@145635.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@145635.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@145635.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@145791.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@145791.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@145791.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@145791.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@145791.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@145791.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@145791.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@145947.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@145947.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@145947.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@145947.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@145947.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@145947.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@145947.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@146103.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@146103.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@146103.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@146103.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@146103.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@146103.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@146103.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@146103.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@144579.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@145485.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@145635.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@145791.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@145947.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@146103.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@145503.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@145499.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@145495.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@145494.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@145493.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@145492.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@145490.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@145489.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@145790.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@145788.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@145787.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@145780.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@145778.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@145776.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@145775.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@145768.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@145766.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@145765.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@145764.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@145763.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@145755.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@145750.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@145946.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@145944.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@145943.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@145936.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@145934.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@145932.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@145931.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@145924.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@145922.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@145921.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@145920.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@145919.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@145911.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@145906.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@146102.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@146100.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@146099.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@146092.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@146090.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@146088.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@146087.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@146080.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@146078.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@146077.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@146076.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@146075.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@146067.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@146062.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@146258.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@146256.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@146255.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@146248.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@146246.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@146244.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@146243.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@146236.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@146234.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@146233.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@146232.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@146231.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@146223.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@146218.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@145513.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@145517.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@145518.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@145519.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@145606.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@145602.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@145597.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@145596.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@145631.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@145630.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@145629.4]
  assign fringeCommon_clock = clock; // @[:@144580.4]
  assign fringeCommon_reset = reset; // @[:@144581.4 FringeZynq.scala 117:22:@145516.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@145507.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@145508.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@145509.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@145510.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@145514.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@145521.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@145520.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@145605.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@145604.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@145603.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@145601.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@145600.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@145599.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@145598.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@145749.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@145742.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@145639.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@145638.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@145905.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@145898.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@145795.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@145794.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@146061.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@146054.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@145951.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@145950.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@146217.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@146210.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@146107.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@146106.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@145634.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@145633.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@145632.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@145486.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@145487.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@145506.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@145505.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@145504.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@145502.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@145501.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@145500.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@145498.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@145497.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@145496.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@145491.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@145488.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@145511.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@145748.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@145747.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@145746.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@145744.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@145743.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@145741.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@145725.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@145726.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@145727.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@145728.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@145729.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@145730.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@145731.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@145732.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@145733.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@145734.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@145735.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@145736.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@145737.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@145738.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@145739.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@145740.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@145661.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@145662.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@145663.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@145664.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@145665.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@145666.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@145667.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@145668.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@145669.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@145670.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@145671.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@145672.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@145673.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@145674.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@145675.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@145676.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@145677.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@145678.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@145679.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@145680.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@145681.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@145682.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@145683.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@145684.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@145685.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@145686.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@145687.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@145688.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@145689.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@145690.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@145691.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@145692.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@145693.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@145694.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@145695.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@145696.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@145697.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@145698.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@145699.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@145700.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@145701.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@145702.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@145703.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@145704.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@145705.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@145706.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@145707.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@145708.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@145709.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@145710.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@145711.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@145712.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@145713.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@145714.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@145715.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@145716.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@145717.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@145718.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@145719.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@145720.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@145721.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@145722.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@145723.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@145724.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@145660.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@145659.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@145640.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@145779.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@145767.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@145762.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@145754.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@145751.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@145904.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@145903.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@145902.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@145900.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@145899.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@145897.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@145881.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@145882.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@145883.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@145884.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@145885.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@145886.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@145887.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@145888.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@145889.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@145890.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@145891.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@145892.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@145893.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@145894.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@145895.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@145896.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@145817.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@145818.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@145819.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@145820.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@145821.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@145822.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@145823.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@145824.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@145825.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@145826.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@145827.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@145828.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@145829.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@145830.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@145831.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@145832.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@145833.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@145834.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@145835.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@145836.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@145837.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@145838.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@145839.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@145840.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@145841.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@145842.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@145843.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@145844.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@145845.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@145846.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@145847.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@145848.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@145849.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@145850.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@145851.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@145852.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@145853.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@145854.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@145855.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@145856.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@145857.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@145858.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@145859.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@145860.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@145861.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@145862.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@145863.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@145864.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@145865.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@145866.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@145867.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@145868.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@145869.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@145870.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@145871.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@145872.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@145873.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@145874.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@145875.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@145876.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@145877.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@145878.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@145879.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@145880.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@145816.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@145815.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@145796.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@145935.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@145923.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@145918.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@145910.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@145907.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@146060.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@146059.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@146058.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@146056.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@146055.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@146053.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@146037.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@146038.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@146039.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@146040.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@146041.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@146042.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@146043.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@146044.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@146045.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@146046.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@146047.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@146048.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@146049.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@146050.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@146051.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@146052.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@145973.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@145974.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@145975.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@145976.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@145977.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@145978.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@145979.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@145980.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@145981.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@145982.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@145983.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@145984.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@145985.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@145986.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@145987.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@145988.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@145989.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@145990.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@145991.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@145992.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@145993.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@145994.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@145995.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@145996.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@145997.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@145998.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@145999.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@146000.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@146001.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@146002.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@146003.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@146004.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@146005.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@146006.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@146007.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@146008.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@146009.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@146010.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@146011.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@146012.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@146013.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@146014.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@146015.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@146016.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@146017.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@146018.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@146019.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@146020.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@146021.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@146022.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@146023.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@146024.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@146025.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@146026.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@146027.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@146028.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@146029.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@146030.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@146031.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@146032.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@146033.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@146034.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@146035.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@146036.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@145972.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@145971.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@145952.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@146091.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@146079.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@146074.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@146066.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@146063.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@146216.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@146215.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@146214.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@146212.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@146211.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@146209.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@146193.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@146194.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@146195.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@146196.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@146197.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@146198.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@146199.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@146200.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@146201.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@146202.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@146203.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@146204.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@146205.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@146206.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@146207.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@146208.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@146129.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@146130.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@146131.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@146132.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@146133.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@146134.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@146135.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@146136.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@146137.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@146138.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@146139.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@146140.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@146141.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@146142.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@146143.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@146144.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@146145.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@146146.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@146147.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@146148.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@146149.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@146150.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@146151.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@146152.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@146153.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@146154.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@146155.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@146156.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@146157.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@146158.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@146159.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@146160.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@146161.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@146162.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@146163.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@146164.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@146165.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@146166.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@146167.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@146168.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@146169.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@146170.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@146171.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@146172.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@146173.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@146174.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@146175.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@146176.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@146177.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@146178.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@146179.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@146180.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@146181.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@146182.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@146183.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@146184.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@146185.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@146186.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@146187.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@146188.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@146189.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@146190.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@146191.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@146192.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@146128.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@146127.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@146108.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@146247.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@146235.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@146230.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@146222.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@146219.4]
endmodule
module SpatialIP( // @[:@146260.2]
  input          clock, // @[:@146261.4]
  input          reset, // @[:@146262.4]
  input          io_raddr, // @[:@146263.4]
  input          io_wen, // @[:@146263.4]
  input          io_waddr, // @[:@146263.4]
  input          io_wdata, // @[:@146263.4]
  output         io_rdata, // @[:@146263.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@146263.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@146263.4]
  input          io_S_AXI_AWVALID, // @[:@146263.4]
  output         io_S_AXI_AWREADY, // @[:@146263.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@146263.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@146263.4]
  input          io_S_AXI_ARVALID, // @[:@146263.4]
  output         io_S_AXI_ARREADY, // @[:@146263.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@146263.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@146263.4]
  input          io_S_AXI_WVALID, // @[:@146263.4]
  output         io_S_AXI_WREADY, // @[:@146263.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@146263.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@146263.4]
  output         io_S_AXI_RVALID, // @[:@146263.4]
  input          io_S_AXI_RREADY, // @[:@146263.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@146263.4]
  output         io_S_AXI_BVALID, // @[:@146263.4]
  input          io_S_AXI_BREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@146263.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@146263.4]
  output         io_M_AXI_0_AWLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@146263.4]
  output         io_M_AXI_0_AWVALID, // @[:@146263.4]
  input          io_M_AXI_0_AWREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@146263.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@146263.4]
  output         io_M_AXI_0_ARLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@146263.4]
  output         io_M_AXI_0_ARVALID, // @[:@146263.4]
  input          io_M_AXI_0_ARREADY, // @[:@146263.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@146263.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@146263.4]
  output         io_M_AXI_0_WLAST, // @[:@146263.4]
  output         io_M_AXI_0_WVALID, // @[:@146263.4]
  input          io_M_AXI_0_WREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@146263.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@146263.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@146263.4]
  input          io_M_AXI_0_RLAST, // @[:@146263.4]
  input          io_M_AXI_0_RVALID, // @[:@146263.4]
  output         io_M_AXI_0_RREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@146263.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@146263.4]
  input          io_M_AXI_0_BVALID, // @[:@146263.4]
  output         io_M_AXI_0_BREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@146263.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@146263.4]
  output         io_M_AXI_1_AWLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@146263.4]
  output         io_M_AXI_1_AWVALID, // @[:@146263.4]
  input          io_M_AXI_1_AWREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@146263.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@146263.4]
  output         io_M_AXI_1_ARLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@146263.4]
  output         io_M_AXI_1_ARVALID, // @[:@146263.4]
  input          io_M_AXI_1_ARREADY, // @[:@146263.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@146263.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@146263.4]
  output         io_M_AXI_1_WLAST, // @[:@146263.4]
  output         io_M_AXI_1_WVALID, // @[:@146263.4]
  input          io_M_AXI_1_WREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@146263.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@146263.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@146263.4]
  input          io_M_AXI_1_RLAST, // @[:@146263.4]
  input          io_M_AXI_1_RVALID, // @[:@146263.4]
  output         io_M_AXI_1_RREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@146263.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@146263.4]
  input          io_M_AXI_1_BVALID, // @[:@146263.4]
  output         io_M_AXI_1_BREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@146263.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@146263.4]
  output         io_M_AXI_2_AWLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@146263.4]
  output         io_M_AXI_2_AWVALID, // @[:@146263.4]
  input          io_M_AXI_2_AWREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@146263.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@146263.4]
  output         io_M_AXI_2_ARLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@146263.4]
  output         io_M_AXI_2_ARVALID, // @[:@146263.4]
  input          io_M_AXI_2_ARREADY, // @[:@146263.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@146263.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@146263.4]
  output         io_M_AXI_2_WLAST, // @[:@146263.4]
  output         io_M_AXI_2_WVALID, // @[:@146263.4]
  input          io_M_AXI_2_WREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@146263.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@146263.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@146263.4]
  input          io_M_AXI_2_RLAST, // @[:@146263.4]
  input          io_M_AXI_2_RVALID, // @[:@146263.4]
  output         io_M_AXI_2_RREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@146263.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@146263.4]
  input          io_M_AXI_2_BVALID, // @[:@146263.4]
  output         io_M_AXI_2_BREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@146263.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@146263.4]
  output         io_M_AXI_3_AWLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@146263.4]
  output         io_M_AXI_3_AWVALID, // @[:@146263.4]
  input          io_M_AXI_3_AWREADY, // @[:@146263.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@146263.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@146263.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@146263.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@146263.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@146263.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@146263.4]
  output         io_M_AXI_3_ARLOCK, // @[:@146263.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@146263.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@146263.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@146263.4]
  output         io_M_AXI_3_ARVALID, // @[:@146263.4]
  input          io_M_AXI_3_ARREADY, // @[:@146263.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@146263.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@146263.4]
  output         io_M_AXI_3_WLAST, // @[:@146263.4]
  output         io_M_AXI_3_WVALID, // @[:@146263.4]
  input          io_M_AXI_3_WREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@146263.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@146263.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@146263.4]
  input          io_M_AXI_3_RLAST, // @[:@146263.4]
  input          io_M_AXI_3_RVALID, // @[:@146263.4]
  output         io_M_AXI_3_RREADY, // @[:@146263.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@146263.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@146263.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@146263.4]
  input          io_M_AXI_3_BVALID, // @[:@146263.4]
  output         io_M_AXI_3_BREADY, // @[:@146263.4]
  input          io_TOP_AXI_AWID, // @[:@146263.4]
  input          io_TOP_AXI_AWUSER, // @[:@146263.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@146263.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@146263.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@146263.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@146263.4]
  input          io_TOP_AXI_AWLOCK, // @[:@146263.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@146263.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@146263.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@146263.4]
  input          io_TOP_AXI_AWVALID, // @[:@146263.4]
  input          io_TOP_AXI_AWREADY, // @[:@146263.4]
  input          io_TOP_AXI_ARID, // @[:@146263.4]
  input          io_TOP_AXI_ARUSER, // @[:@146263.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@146263.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@146263.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@146263.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@146263.4]
  input          io_TOP_AXI_ARLOCK, // @[:@146263.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@146263.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@146263.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@146263.4]
  input          io_TOP_AXI_ARVALID, // @[:@146263.4]
  input          io_TOP_AXI_ARREADY, // @[:@146263.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@146263.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@146263.4]
  input          io_TOP_AXI_WLAST, // @[:@146263.4]
  input          io_TOP_AXI_WVALID, // @[:@146263.4]
  input          io_TOP_AXI_WREADY, // @[:@146263.4]
  input          io_TOP_AXI_RID, // @[:@146263.4]
  input          io_TOP_AXI_RUSER, // @[:@146263.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@146263.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@146263.4]
  input          io_TOP_AXI_RLAST, // @[:@146263.4]
  input          io_TOP_AXI_RVALID, // @[:@146263.4]
  input          io_TOP_AXI_RREADY, // @[:@146263.4]
  input          io_TOP_AXI_BID, // @[:@146263.4]
  input          io_TOP_AXI_BUSER, // @[:@146263.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@146263.4]
  input          io_TOP_AXI_BVALID, // @[:@146263.4]
  input          io_TOP_AXI_BREADY, // @[:@146263.4]
  input          io_DWIDTH_AXI_AWID, // @[:@146263.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@146263.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@146263.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@146263.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@146263.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@146263.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@146263.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@146263.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@146263.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@146263.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@146263.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@146263.4]
  input          io_DWIDTH_AXI_ARID, // @[:@146263.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@146263.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@146263.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@146263.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@146263.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@146263.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@146263.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@146263.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@146263.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@146263.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@146263.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@146263.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@146263.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@146263.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@146263.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@146263.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@146263.4]
  input          io_DWIDTH_AXI_RID, // @[:@146263.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@146263.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@146263.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@146263.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@146263.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@146263.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@146263.4]
  input          io_DWIDTH_AXI_BID, // @[:@146263.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@146263.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@146263.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@146263.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@146263.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@146263.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@146263.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@146263.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@146263.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@146263.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@146263.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@146263.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@146263.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@146263.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@146263.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@146263.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@146263.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@146263.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@146263.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@146263.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@146263.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@146263.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@146263.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@146263.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@146263.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@146263.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@146263.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@146263.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@146263.4]
  input          io_PROTOCOL_AXI_RID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@146263.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@146263.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@146263.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@146263.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@146263.4]
  input          io_PROTOCOL_AXI_BID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@146263.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@146263.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@146263.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@146263.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@146263.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@146263.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@146263.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@146263.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@146263.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@146263.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@146263.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@146263.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@146263.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@146263.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@146263.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@146263.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@146263.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@146263.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@146263.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@146263.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@146263.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@146263.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@146263.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@146263.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@146265.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@146265.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@146265.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@146265.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@146265.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@146265.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@146265.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@146265.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@146265.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@146265.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@146407.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@146407.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@146407.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@146407.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@146407.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@146407.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@146407.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@146265.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@146407.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@146425.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@146421.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@146417.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@146416.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@146415.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@146414.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@146412.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@146411.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@146469.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146468.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@146467.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@146466.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146465.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146464.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146463.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146462.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146461.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146460.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@146459.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@146457.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146456.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@146455.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@146454.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146453.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146452.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146451.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146450.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146449.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146448.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@146447.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@146445.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@146444.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@146443.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@146442.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@146434.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@146429.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@146510.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146509.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@146508.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@146507.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146506.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146505.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146504.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146503.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146502.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146501.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@146500.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@146498.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146497.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@146496.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@146495.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146494.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146493.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146492.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146491.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146490.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146489.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@146488.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@146486.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@146485.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@146484.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@146483.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@146475.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@146470.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@146551.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146550.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@146549.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@146548.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146547.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146546.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146545.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146544.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146543.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146542.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@146541.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@146539.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146538.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@146537.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@146536.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146535.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146534.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146533.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146532.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146531.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146530.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@146529.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@146527.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@146526.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@146525.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@146524.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@146516.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@146511.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@146592.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146591.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@146590.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@146589.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146588.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146587.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146586.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146585.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146584.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146583.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@146582.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@146580.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146579.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@146578.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@146577.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146576.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146575.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146574.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146573.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146572.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146571.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@146570.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@146568.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@146567.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@146566.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@146565.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@146557.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@146552.4]
  assign accel_clock = clock; // @[:@146266.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@146267.4 Zynq.scala 54:17:@146881.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@146876.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@146869.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@146864.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@146848.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@146849.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@146850.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@146851.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@146852.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@146853.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@146854.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@146855.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@146856.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@146857.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@146858.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@146859.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@146860.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@146861.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@146862.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@146863.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@146847.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@146843.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@146838.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@146837.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@146836.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@146817.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@146801.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@146802.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@146803.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@146804.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@146805.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@146806.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@146807.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@146808.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@146809.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@146810.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@146811.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@146812.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@146813.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@146814.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@146815.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@146816.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@146800.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@146765.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@146764.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@146872.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@146871.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@146870.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@146758.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@146759.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@146762.4]
  assign FringeZynq_clock = clock; // @[:@146408.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@146409.4 Zynq.scala 53:18:@146880.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@146428.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@146427.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@146426.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@146424.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@146423.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@146422.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@146420.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@146419.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@146418.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@146413.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@146410.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@146458.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@146446.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@146441.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@146433.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@146430.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@146499.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@146487.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@146482.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@146474.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@146471.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@146540.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@146528.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@146523.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@146515.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@146512.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@146581.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@146569.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@146564.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@146556.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@146553.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@146877.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@146761.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@146760.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@146846.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@146845.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@146844.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@146842.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@146841.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@146840.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@146839.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@146875.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@146874.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@146873.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




