module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  output [31:0] O_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x201_TREADY(dontcare), // @[:@1298.4]
    .io_in_x201_TDATA(I_0), // @[:@1298.4]
    .io_in_x201_TID(8'h0),
    .io_in_x201_TDEST(8'h0),
    .io_in_x202_TVALID(valid_down), // @[:@1298.4]
    .io_in_x202_TDATA(O_0), // @[:@1298.4]
    .io_in_x202_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x209_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(reset), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule

module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh54); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh54); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x203_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x491_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x359_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x204_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x205_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x209_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x222_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x408_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x215_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x222_inr_Foreach_kernelx222_inr_Foreach_concrete1( // @[:@4533.2]
  input         clock, // @[:@4534.4]
  input         reset, // @[:@4535.4]
  output        io_in_x205_fifoinpacked_0_wPort_0_en_0, // @[:@4536.4]
  input         io_in_x205_fifoinpacked_0_full, // @[:@4536.4]
  output        io_in_x205_fifoinpacked_0_active_0_in, // @[:@4536.4]
  input         io_in_x205_fifoinpacked_0_active_0_out, // @[:@4536.4]
  input         io_sigsIn_backpressure, // @[:@4536.4]
  input         io_sigsIn_datapathEn, // @[:@4536.4]
  input         io_sigsIn_break, // @[:@4536.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@4536.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4536.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4536.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@4536.4]
  input         io_rr // @[:@4536.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4570.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4570.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4582.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@4582.4]
  wire  x408_sub_1_clock; // @[Math.scala 191:24:@4609.4]
  wire  x408_sub_1_reset; // @[Math.scala 191:24:@4609.4]
  wire [31:0] x408_sub_1_io_a; // @[Math.scala 191:24:@4609.4]
  wire [31:0] x408_sub_1_io_b; // @[Math.scala 191:24:@4609.4]
  wire  x408_sub_1_io_flow; // @[Math.scala 191:24:@4609.4]
  wire [31:0] x408_sub_1_io_result; // @[Math.scala 191:24:@4609.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4619.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4619.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4619.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4619.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4619.4]
  wire  x215_sum_1_clock; // @[Math.scala 150:24:@4628.4]
  wire  x215_sum_1_reset; // @[Math.scala 150:24:@4628.4]
  wire [31:0] x215_sum_1_io_a; // @[Math.scala 150:24:@4628.4]
  wire [31:0] x215_sum_1_io_b; // @[Math.scala 150:24:@4628.4]
  wire  x215_sum_1_io_flow; // @[Math.scala 150:24:@4628.4]
  wire [31:0] x215_sum_1_io_result; // @[Math.scala 150:24:@4628.4]
  wire  x216_sum_1_clock; // @[Math.scala 150:24:@4640.4]
  wire  x216_sum_1_reset; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x216_sum_1_io_a; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x216_sum_1_io_b; // @[Math.scala 150:24:@4640.4]
  wire  x216_sum_1_io_flow; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x216_sum_1_io_result; // @[Math.scala 150:24:@4640.4]
  wire [31:0] x218_1_io_b; // @[Math.scala 720:24:@4661.4]
  wire [31:0] x218_1_io_result; // @[Math.scala 720:24:@4661.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4674.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4683.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4694.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4694.4]
  wire  _T_327; // @[sm_x222_inr_Foreach.scala 62:18:@4595.4]
  wire  _T_328; // @[sm_x222_inr_Foreach.scala 62:55:@4596.4]
  wire [31:0] b210_number; // @[Math.scala 723:22:@4575.4 Math.scala 724:14:@4576.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@4600.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@4600.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@4605.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@4605.4]
  wire [31:0] x216_sum_number; // @[Math.scala 154:22:@4646.4 Math.scala 155:14:@4647.4]
  wire [31:0] _T_358; // @[Math.scala 406:49:@4653.4]
  wire [31:0] _T_360; // @[Math.scala 406:56:@4655.4]
  wire [31:0] _T_361; // @[Math.scala 406:56:@4656.4]
  wire  _T_379; // @[sm_x222_inr_Foreach.scala 89:131:@4691.4]
  wire  _T_383; // @[package.scala 96:25:@4699.4 package.scala 96:25:@4700.4]
  wire  _T_385; // @[implicits.scala 55:10:@4701.4]
  wire  _T_386; // @[sm_x222_inr_Foreach.scala 89:148:@4702.4]
  wire  _T_388; // @[sm_x222_inr_Foreach.scala 89:236:@4704.4]
  wire  _T_389; // @[sm_x222_inr_Foreach.scala 89:255:@4705.4]
  wire  x495_b212_D3; // @[package.scala 96:25:@4688.4 package.scala 96:25:@4689.4]
  wire  _T_392; // @[sm_x222_inr_Foreach.scala 89:291:@4707.4]
  wire  x494_b213_D3; // @[package.scala 96:25:@4679.4 package.scala 96:25:@4680.4]
  _ _ ( // @[Math.scala 720:24:@4570.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@4582.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x408_sub x408_sub_1 ( // @[Math.scala 191:24:@4609.4]
    .clock(x408_sub_1_clock),
    .reset(x408_sub_1_reset),
    .io_a(x408_sub_1_io_a),
    .io_b(x408_sub_1_io_b),
    .io_flow(x408_sub_1_io_flow),
    .io_result(x408_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@4619.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x215_sum x215_sum_1 ( // @[Math.scala 150:24:@4628.4]
    .clock(x215_sum_1_clock),
    .reset(x215_sum_1_reset),
    .io_a(x215_sum_1_io_a),
    .io_b(x215_sum_1_io_b),
    .io_flow(x215_sum_1_io_flow),
    .io_result(x215_sum_1_io_result)
  );
  x215_sum x216_sum_1 ( // @[Math.scala 150:24:@4640.4]
    .clock(x216_sum_1_clock),
    .reset(x216_sum_1_reset),
    .io_a(x216_sum_1_io_a),
    .io_b(x216_sum_1_io_b),
    .io_flow(x216_sum_1_io_flow),
    .io_result(x216_sum_1_io_result)
  );
  _ x218_1 ( // @[Math.scala 720:24:@4661.4]
    .io_b(x218_1_io_b),
    .io_result(x218_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4674.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@4683.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@4694.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x205_fifoinpacked_0_full; // @[sm_x222_inr_Foreach.scala 62:18:@4595.4]
  assign _T_328 = ~ io_in_x205_fifoinpacked_0_active_0_out; // @[sm_x222_inr_Foreach.scala 62:55:@4596.4]
  assign b210_number = __io_result; // @[Math.scala 723:22:@4575.4 Math.scala 724:14:@4576.4]
  assign _GEN_0 = {{11'd0}, b210_number}; // @[Math.scala 461:32:@4600.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@4600.4]
  assign _GEN_1 = {{7'd0}, b210_number}; // @[Math.scala 461:32:@4605.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@4605.4]
  assign x216_sum_number = x216_sum_1_io_result; // @[Math.scala 154:22:@4646.4 Math.scala 155:14:@4647.4]
  assign _T_358 = $signed(x216_sum_number); // @[Math.scala 406:49:@4653.4]
  assign _T_360 = $signed(_T_358) & $signed(32'shff); // @[Math.scala 406:56:@4655.4]
  assign _T_361 = $signed(_T_360); // @[Math.scala 406:56:@4656.4]
  assign _T_379 = ~ io_sigsIn_break; // @[sm_x222_inr_Foreach.scala 89:131:@4691.4]
  assign _T_383 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4699.4 package.scala 96:25:@4700.4]
  assign _T_385 = io_rr ? _T_383 : 1'h0; // @[implicits.scala 55:10:@4701.4]
  assign _T_386 = _T_379 & _T_385; // @[sm_x222_inr_Foreach.scala 89:148:@4702.4]
  assign _T_388 = _T_386 & _T_379; // @[sm_x222_inr_Foreach.scala 89:236:@4704.4]
  assign _T_389 = _T_388 & io_sigsIn_backpressure; // @[sm_x222_inr_Foreach.scala 89:255:@4705.4]
  assign x495_b212_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4688.4 package.scala 96:25:@4689.4]
  assign _T_392 = _T_389 & x495_b212_D3; // @[sm_x222_inr_Foreach.scala 89:291:@4707.4]
  assign x494_b213_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4679.4 package.scala 96:25:@4680.4]
  assign io_in_x205_fifoinpacked_0_wPort_0_en_0 = _T_392 & x494_b213_D3; // @[MemInterfaceType.scala 93:57:@4711.4]
  assign io_in_x205_fifoinpacked_0_active_0_in = x495_b212_D3 & x494_b213_D3; // @[MemInterfaceType.scala 147:18:@4714.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4573.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@4585.4]
  assign x408_sub_1_clock = clock; // @[:@4610.4]
  assign x408_sub_1_reset = reset; // @[:@4611.4]
  assign x408_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@4612.4]
  assign x408_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@4613.4]
  assign x408_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@4614.4]
  assign RetimeWrapper_clock = clock; // @[:@4620.4]
  assign RetimeWrapper_reset = reset; // @[:@4621.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4623.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@4622.4]
  assign x215_sum_1_clock = clock; // @[:@4629.4]
  assign x215_sum_1_reset = reset; // @[:@4630.4]
  assign x215_sum_1_io_a = x408_sub_1_io_result; // @[Math.scala 151:17:@4631.4]
  assign x215_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@4632.4]
  assign x215_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4633.4]
  assign x216_sum_1_clock = clock; // @[:@4641.4]
  assign x216_sum_1_reset = reset; // @[:@4642.4]
  assign x216_sum_1_io_a = x215_sum_1_io_result; // @[Math.scala 151:17:@4643.4]
  assign x216_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@4644.4]
  assign x216_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4645.4]
  assign x218_1_io_b = $unsigned(_T_361); // @[Math.scala 721:17:@4664.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4675.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4676.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4678.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@4677.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4684.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4685.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4687.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4686.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4695.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4696.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4698.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4697.4]
endmodule
module RetimeWrapper_41( // @[:@5832.2]
  input   clock, // @[:@5833.4]
  input   reset, // @[:@5834.4]
  input   io_flow, // @[:@5835.4]
  input   io_in, // @[:@5835.4]
  output  io_out // @[:@5835.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5837.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(169)) sr ( // @[RetimeShiftRegister.scala 15:20:@5837.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5850.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5849.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5848.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5847.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5846.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5844.4]
endmodule
module RetimeWrapper_45( // @[:@5960.2]
  input   clock, // @[:@5961.4]
  input   reset, // @[:@5962.4]
  input   io_flow, // @[:@5963.4]
  input   io_in, // @[:@5963.4]
  output  io_out // @[:@5963.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5965.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(168)) sr ( // @[RetimeShiftRegister.scala 15:20:@5965.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5978.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5977.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5976.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5975.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5974.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5972.4]
endmodule
module x357_inr_Foreach_SAMPLER_BOX_sm( // @[:@5980.2]
  input   clock, // @[:@5981.4]
  input   reset, // @[:@5982.4]
  input   io_enable, // @[:@5983.4]
  output  io_done, // @[:@5983.4]
  output  io_doneLatch, // @[:@5983.4]
  input   io_ctrDone, // @[:@5983.4]
  output  io_datapathEn, // @[:@5983.4]
  output  io_ctrInc, // @[:@5983.4]
  output  io_ctrRst, // @[:@5983.4]
  input   io_parentAck, // @[:@5983.4]
  input   io_backpressure, // @[:@5983.4]
  input   io_break // @[:@5983.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@5985.4]
  wire  active_reset; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@5985.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@5985.4]
  wire  done_clock; // @[Controllers.scala 262:20:@5988.4]
  wire  done_reset; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@5988.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@5988.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6022.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6044.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6056.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6064.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6080.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6080.4]
  wire  _T_80; // @[Controllers.scala 264:48:@5993.4]
  wire  _T_81; // @[Controllers.scala 264:46:@5994.4]
  wire  _T_82; // @[Controllers.scala 264:62:@5995.4]
  wire  _T_83; // @[Controllers.scala 264:60:@5996.4]
  wire  _T_100; // @[package.scala 100:49:@6013.4]
  reg  _T_103; // @[package.scala 48:56:@6014.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6027.4 package.scala 96:25:@6028.4]
  wire  _T_110; // @[package.scala 100:49:@6029.4]
  reg  _T_113; // @[package.scala 48:56:@6030.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6032.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6037.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6038.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6041.4]
  wire  _T_124; // @[package.scala 96:25:@6049.4 package.scala 96:25:@6050.4]
  wire  _T_126; // @[package.scala 100:49:@6051.4]
  reg  _T_129; // @[package.scala 48:56:@6052.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6074.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6076.4]
  reg  _T_153; // @[package.scala 48:56:@6077.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6085.4 package.scala 96:25:@6086.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6087.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6088.4]
  SRFF active ( // @[Controllers.scala 261:22:@5985.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@5988.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_41 RetimeWrapper ( // @[package.scala 93:22:@6022.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_41 RetimeWrapper_1 ( // @[package.scala 93:22:@6044.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6056.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6064.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_45 RetimeWrapper_4 ( // @[package.scala 93:22:@6080.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@5993.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@5994.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@5995.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@5996.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6013.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6027.4 package.scala 96:25:@6028.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6029.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6032.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6037.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6038.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6041.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6049.4 package.scala 96:25:@6050.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6051.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6076.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6085.4 package.scala 96:25:@6086.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6087.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6088.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6055.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6090.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6040.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6043.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6035.4]
  assign active_clock = clock; // @[:@5986.4]
  assign active_reset = reset; // @[:@5987.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@5998.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6002.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6003.4]
  assign done_clock = clock; // @[:@5989.4]
  assign done_reset = reset; // @[:@5990.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6018.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6011.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6012.4]
  assign RetimeWrapper_clock = clock; // @[:@6023.4]
  assign RetimeWrapper_reset = reset; // @[:@6024.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6026.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6025.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6045.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6046.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6048.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6047.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6057.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6058.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6060.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6059.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6065.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6066.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6068.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6067.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6081.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6082.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6084.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6083.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SRAM_1( // @[:@6317.2]
  input         clock, // @[:@6318.4]
  input         reset, // @[:@6319.4]
  input  [9:0]  io_raddr, // @[:@6320.4]
  input         io_wen, // @[:@6320.4]
  input  [9:0]  io_waddr, // @[:@6320.4]
  input  [31:0] io_wdata, // @[:@6320.4]
  output [31:0] io_rdata, // @[:@6320.4]
  input         io_backpressure // @[:@6320.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6322.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6322.4]
  wire [9:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6322.4]
  wire [9:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6322.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6322.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6340.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6341.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6342.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6344.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(640), .AWIDTH(10)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6322.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6340.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6341.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6349.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6336.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6337.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6334.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6339.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6338.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6335.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6333.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6332.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_50( // @[:@6363.2]
  input        clock, // @[:@6364.4]
  input        reset, // @[:@6365.4]
  input        io_flow, // @[:@6366.4]
  input  [9:0] io_in, // @[:@6366.4]
  output [9:0] io_out // @[:@6366.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6368.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6368.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6381.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6380.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@6379.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6378.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6377.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6375.4]
endmodule
module Mem1D_5( // @[:@6383.2]
  input         clock, // @[:@6384.4]
  input         reset, // @[:@6385.4]
  input  [9:0]  io_r_ofs_0, // @[:@6386.4]
  input         io_r_backpressure, // @[:@6386.4]
  input  [9:0]  io_w_ofs_0, // @[:@6386.4]
  input  [31:0] io_w_data_0, // @[:@6386.4]
  input         io_w_en_0, // @[:@6386.4]
  output [31:0] io_output // @[:@6386.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [9:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [9:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@6390.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@6390.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6393.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6393.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6393.4]
  wire [9:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6393.4]
  wire [9:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6393.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@6388.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@6390.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@6393.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 10'h280; // @[MemPrimitives.scala 702:32:@6388.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@6406.4]
  assign SRAM_clock = clock; // @[:@6391.4]
  assign SRAM_reset = reset; // @[:@6392.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@6400.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@6403.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@6401.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@6404.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@6405.4]
  assign RetimeWrapper_clock = clock; // @[:@6394.4]
  assign RetimeWrapper_reset = reset; // @[:@6395.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@6397.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@6396.4]
endmodule
module StickySelects_1( // @[:@7585.2]
  input   clock, // @[:@7586.4]
  input   reset, // @[:@7587.4]
  input   io_ins_0, // @[:@7588.4]
  input   io_ins_1, // @[:@7588.4]
  input   io_ins_2, // @[:@7588.4]
  input   io_ins_3, // @[:@7588.4]
  input   io_ins_4, // @[:@7588.4]
  input   io_ins_5, // @[:@7588.4]
  input   io_ins_6, // @[:@7588.4]
  input   io_ins_7, // @[:@7588.4]
  input   io_ins_8, // @[:@7588.4]
  output  io_outs_0, // @[:@7588.4]
  output  io_outs_1, // @[:@7588.4]
  output  io_outs_2, // @[:@7588.4]
  output  io_outs_3, // @[:@7588.4]
  output  io_outs_4, // @[:@7588.4]
  output  io_outs_5, // @[:@7588.4]
  output  io_outs_6, // @[:@7588.4]
  output  io_outs_7, // @[:@7588.4]
  output  io_outs_8 // @[:@7588.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@7590.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@7591.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@7592.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@7593.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@7594.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@7595.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@7596.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@7597.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@7598.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@7599.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@7600.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@7601.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@7602.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@7603.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@7604.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@7605.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@7606.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@7607.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@7609.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@7610.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@7611.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@7612.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@7613.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@7614.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@7615.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@7616.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@7617.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@7619.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@7620.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@7621.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@7622.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@7623.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@7624.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@7625.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@7626.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@7627.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@7630.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@7631.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@7632.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@7633.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@7634.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@7635.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@7636.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@7637.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@7641.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@7642.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@7643.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@7644.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@7645.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@7646.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@7647.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@7652.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@7653.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@7654.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@7655.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@7656.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@7657.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@7663.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@7664.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@7665.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@7666.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@7667.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@7674.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@7675.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@7676.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@7677.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@7685.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@7686.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@7687.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@7599.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@7600.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@7601.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@7602.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@7603.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@7604.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@7605.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@7606.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@7607.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@7609.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@7610.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@7611.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@7612.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@7613.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@7614.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@7615.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@7616.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@7617.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@7619.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@7620.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@7621.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@7622.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@7623.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@7624.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@7625.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@7626.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@7627.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@7630.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@7631.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@7632.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@7633.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@7634.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@7635.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@7636.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@7637.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@7641.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@7642.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@7643.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@7644.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@7645.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@7646.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@7647.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@7652.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@7653.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@7654.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@7655.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@7656.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@7657.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@7663.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@7664.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@7665.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@7666.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@7667.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@7674.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@7675.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@7676.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@7677.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@7685.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@7686.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@7687.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@7689.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@7690.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@7691.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@7692.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@7693.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@7694.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@7695.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@7696.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@7697.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x233_lb_0( // @[:@12409.2]
  input         clock, // @[:@12410.4]
  input         reset, // @[:@12411.4]
  input  [1:0]  io_rPort_8_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_8_ofs_0, // @[:@12412.4]
  input         io_rPort_8_en_0, // @[:@12412.4]
  input         io_rPort_8_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_8_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_7_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_7_ofs_0, // @[:@12412.4]
  input         io_rPort_7_en_0, // @[:@12412.4]
  input         io_rPort_7_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_7_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_6_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_6_ofs_0, // @[:@12412.4]
  input         io_rPort_6_en_0, // @[:@12412.4]
  input         io_rPort_6_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_6_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_5_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_5_ofs_0, // @[:@12412.4]
  input         io_rPort_5_en_0, // @[:@12412.4]
  input         io_rPort_5_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_5_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_4_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_4_ofs_0, // @[:@12412.4]
  input         io_rPort_4_en_0, // @[:@12412.4]
  input         io_rPort_4_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_4_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_3_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_3_ofs_0, // @[:@12412.4]
  input         io_rPort_3_en_0, // @[:@12412.4]
  input         io_rPort_3_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_3_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_2_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_2_ofs_0, // @[:@12412.4]
  input         io_rPort_2_en_0, // @[:@12412.4]
  input         io_rPort_2_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_2_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_1_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_1_ofs_0, // @[:@12412.4]
  input         io_rPort_1_en_0, // @[:@12412.4]
  input         io_rPort_1_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_1_output_0, // @[:@12412.4]
  input  [1:0]  io_rPort_0_banks_1, // @[:@12412.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12412.4]
  input  [9:0]  io_rPort_0_ofs_0, // @[:@12412.4]
  input         io_rPort_0_en_0, // @[:@12412.4]
  input         io_rPort_0_backpressure, // @[:@12412.4]
  output [31:0] io_rPort_0_output_0, // @[:@12412.4]
  input  [1:0]  io_wPort_0_banks_1, // @[:@12412.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12412.4]
  input  [9:0]  io_wPort_0_ofs_0, // @[:@12412.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12412.4]
  input         io_wPort_0_en_0 // @[:@12412.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [9:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [9:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12477.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12477.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [9:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [9:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12493.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12493.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [9:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [9:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12509.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12509.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [9:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [9:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12525.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12525.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [9:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [9:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12541.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12541.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [9:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [9:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12557.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12557.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [9:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [9:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12573.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12573.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [9:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [9:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12589.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12589.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [9:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [9:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12605.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12605.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [9:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [9:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12621.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12621.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [9:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [9:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12637.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12637.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [9:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [9:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12653.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12653.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 124:33:@12849.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 124:33:@12938.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 124:33:@13027.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 124:33:@13116.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 124:33:@13205.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 124:33:@13383.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 124:33:@13472.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 124:33:@13561.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 124:33:@13650.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 124:33:@13739.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 124:33:@13828.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@13918.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@13926.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@13934.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@13942.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@13950.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@13958.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@13966.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@13974.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@13982.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@13990.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@13998.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14006.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14062.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14070.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14078.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14206.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14214.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14222.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14350.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14358.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14366.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14494.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14502.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14510.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14638.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14646.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14654.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14782.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14790.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@14926.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@14942.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@15070.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@15078.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@15086.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@15158.4]
  wire  _T_316; // @[MemPrimitives.scala 82:210:@12669.4]
  wire  _T_318; // @[MemPrimitives.scala 82:210:@12670.4]
  wire  _T_319; // @[MemPrimitives.scala 82:228:@12671.4]
  wire  _T_320; // @[MemPrimitives.scala 83:102:@12672.4]
  wire [42:0] _T_322; // @[Cat.scala 30:58:@12674.4]
  wire  _T_329; // @[MemPrimitives.scala 82:210:@12682.4]
  wire  _T_330; // @[MemPrimitives.scala 82:228:@12683.4]
  wire  _T_331; // @[MemPrimitives.scala 83:102:@12684.4]
  wire [42:0] _T_333; // @[Cat.scala 30:58:@12686.4]
  wire  _T_340; // @[MemPrimitives.scala 82:210:@12694.4]
  wire  _T_341; // @[MemPrimitives.scala 82:228:@12695.4]
  wire  _T_342; // @[MemPrimitives.scala 83:102:@12696.4]
  wire [42:0] _T_344; // @[Cat.scala 30:58:@12698.4]
  wire  _T_349; // @[MemPrimitives.scala 82:210:@12705.4]
  wire  _T_352; // @[MemPrimitives.scala 82:228:@12707.4]
  wire  _T_353; // @[MemPrimitives.scala 83:102:@12708.4]
  wire [42:0] _T_355; // @[Cat.scala 30:58:@12710.4]
  wire  _T_363; // @[MemPrimitives.scala 82:228:@12719.4]
  wire  _T_364; // @[MemPrimitives.scala 83:102:@12720.4]
  wire [42:0] _T_366; // @[Cat.scala 30:58:@12722.4]
  wire  _T_374; // @[MemPrimitives.scala 82:228:@12731.4]
  wire  _T_375; // @[MemPrimitives.scala 83:102:@12732.4]
  wire [42:0] _T_377; // @[Cat.scala 30:58:@12734.4]
  wire  _T_382; // @[MemPrimitives.scala 82:210:@12741.4]
  wire  _T_385; // @[MemPrimitives.scala 82:228:@12743.4]
  wire  _T_386; // @[MemPrimitives.scala 83:102:@12744.4]
  wire [42:0] _T_388; // @[Cat.scala 30:58:@12746.4]
  wire  _T_396; // @[MemPrimitives.scala 82:228:@12755.4]
  wire  _T_397; // @[MemPrimitives.scala 83:102:@12756.4]
  wire [42:0] _T_399; // @[Cat.scala 30:58:@12758.4]
  wire  _T_407; // @[MemPrimitives.scala 82:228:@12767.4]
  wire  _T_408; // @[MemPrimitives.scala 83:102:@12768.4]
  wire [42:0] _T_410; // @[Cat.scala 30:58:@12770.4]
  wire  _T_415; // @[MemPrimitives.scala 82:210:@12777.4]
  wire  _T_418; // @[MemPrimitives.scala 82:228:@12779.4]
  wire  _T_419; // @[MemPrimitives.scala 83:102:@12780.4]
  wire [42:0] _T_421; // @[Cat.scala 30:58:@12782.4]
  wire  _T_429; // @[MemPrimitives.scala 82:228:@12791.4]
  wire  _T_430; // @[MemPrimitives.scala 83:102:@12792.4]
  wire [42:0] _T_432; // @[Cat.scala 30:58:@12794.4]
  wire  _T_440; // @[MemPrimitives.scala 82:228:@12803.4]
  wire  _T_441; // @[MemPrimitives.scala 83:102:@12804.4]
  wire [42:0] _T_443; // @[Cat.scala 30:58:@12806.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@12813.4]
  wire  _T_450; // @[MemPrimitives.scala 110:210:@12814.4]
  wire  _T_451; // @[MemPrimitives.scala 110:228:@12815.4]
  wire  _T_454; // @[MemPrimitives.scala 110:210:@12817.4]
  wire  _T_456; // @[MemPrimitives.scala 110:210:@12818.4]
  wire  _T_457; // @[MemPrimitives.scala 110:228:@12819.4]
  wire  _T_460; // @[MemPrimitives.scala 110:210:@12821.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@12822.4]
  wire  _T_463; // @[MemPrimitives.scala 110:228:@12823.4]
  wire  _T_466; // @[MemPrimitives.scala 110:210:@12825.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@12826.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@12827.4]
  wire  _T_472; // @[MemPrimitives.scala 110:210:@12829.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@12830.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@12831.4]
  wire  _T_478; // @[MemPrimitives.scala 110:210:@12833.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@12834.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@12835.4]
  wire  _T_484; // @[MemPrimitives.scala 110:210:@12837.4]
  wire  _T_486; // @[MemPrimitives.scala 110:210:@12838.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@12839.4]
  wire  _T_490; // @[MemPrimitives.scala 110:210:@12841.4]
  wire  _T_492; // @[MemPrimitives.scala 110:210:@12842.4]
  wire  _T_493; // @[MemPrimitives.scala 110:228:@12843.4]
  wire  _T_496; // @[MemPrimitives.scala 110:210:@12845.4]
  wire  _T_498; // @[MemPrimitives.scala 110:210:@12846.4]
  wire  _T_499; // @[MemPrimitives.scala 110:228:@12847.4]
  wire  _T_501; // @[MemPrimitives.scala 126:35:@12861.4]
  wire  _T_502; // @[MemPrimitives.scala 126:35:@12862.4]
  wire  _T_503; // @[MemPrimitives.scala 126:35:@12863.4]
  wire  _T_504; // @[MemPrimitives.scala 126:35:@12864.4]
  wire  _T_505; // @[MemPrimitives.scala 126:35:@12865.4]
  wire  _T_506; // @[MemPrimitives.scala 126:35:@12866.4]
  wire  _T_507; // @[MemPrimitives.scala 126:35:@12867.4]
  wire  _T_508; // @[MemPrimitives.scala 126:35:@12868.4]
  wire  _T_509; // @[MemPrimitives.scala 126:35:@12869.4]
  wire [11:0] _T_511; // @[Cat.scala 30:58:@12871.4]
  wire [11:0] _T_513; // @[Cat.scala 30:58:@12873.4]
  wire [11:0] _T_515; // @[Cat.scala 30:58:@12875.4]
  wire [11:0] _T_517; // @[Cat.scala 30:58:@12877.4]
  wire [11:0] _T_519; // @[Cat.scala 30:58:@12879.4]
  wire [11:0] _T_521; // @[Cat.scala 30:58:@12881.4]
  wire [11:0] _T_523; // @[Cat.scala 30:58:@12883.4]
  wire [11:0] _T_525; // @[Cat.scala 30:58:@12885.4]
  wire [11:0] _T_527; // @[Cat.scala 30:58:@12887.4]
  wire [11:0] _T_528; // @[Mux.scala 31:69:@12888.4]
  wire [11:0] _T_529; // @[Mux.scala 31:69:@12889.4]
  wire [11:0] _T_530; // @[Mux.scala 31:69:@12890.4]
  wire [11:0] _T_531; // @[Mux.scala 31:69:@12891.4]
  wire [11:0] _T_532; // @[Mux.scala 31:69:@12892.4]
  wire [11:0] _T_533; // @[Mux.scala 31:69:@12893.4]
  wire [11:0] _T_534; // @[Mux.scala 31:69:@12894.4]
  wire [11:0] _T_535; // @[Mux.scala 31:69:@12895.4]
  wire  _T_542; // @[MemPrimitives.scala 110:210:@12903.4]
  wire  _T_543; // @[MemPrimitives.scala 110:228:@12904.4]
  wire  _T_548; // @[MemPrimitives.scala 110:210:@12907.4]
  wire  _T_549; // @[MemPrimitives.scala 110:228:@12908.4]
  wire  _T_554; // @[MemPrimitives.scala 110:210:@12911.4]
  wire  _T_555; // @[MemPrimitives.scala 110:228:@12912.4]
  wire  _T_560; // @[MemPrimitives.scala 110:210:@12915.4]
  wire  _T_561; // @[MemPrimitives.scala 110:228:@12916.4]
  wire  _T_566; // @[MemPrimitives.scala 110:210:@12919.4]
  wire  _T_567; // @[MemPrimitives.scala 110:228:@12920.4]
  wire  _T_572; // @[MemPrimitives.scala 110:210:@12923.4]
  wire  _T_573; // @[MemPrimitives.scala 110:228:@12924.4]
  wire  _T_578; // @[MemPrimitives.scala 110:210:@12927.4]
  wire  _T_579; // @[MemPrimitives.scala 110:228:@12928.4]
  wire  _T_584; // @[MemPrimitives.scala 110:210:@12931.4]
  wire  _T_585; // @[MemPrimitives.scala 110:228:@12932.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@12935.4]
  wire  _T_591; // @[MemPrimitives.scala 110:228:@12936.4]
  wire  _T_593; // @[MemPrimitives.scala 126:35:@12950.4]
  wire  _T_594; // @[MemPrimitives.scala 126:35:@12951.4]
  wire  _T_595; // @[MemPrimitives.scala 126:35:@12952.4]
  wire  _T_596; // @[MemPrimitives.scala 126:35:@12953.4]
  wire  _T_597; // @[MemPrimitives.scala 126:35:@12954.4]
  wire  _T_598; // @[MemPrimitives.scala 126:35:@12955.4]
  wire  _T_599; // @[MemPrimitives.scala 126:35:@12956.4]
  wire  _T_600; // @[MemPrimitives.scala 126:35:@12957.4]
  wire  _T_601; // @[MemPrimitives.scala 126:35:@12958.4]
  wire [11:0] _T_603; // @[Cat.scala 30:58:@12960.4]
  wire [11:0] _T_605; // @[Cat.scala 30:58:@12962.4]
  wire [11:0] _T_607; // @[Cat.scala 30:58:@12964.4]
  wire [11:0] _T_609; // @[Cat.scala 30:58:@12966.4]
  wire [11:0] _T_611; // @[Cat.scala 30:58:@12968.4]
  wire [11:0] _T_613; // @[Cat.scala 30:58:@12970.4]
  wire [11:0] _T_615; // @[Cat.scala 30:58:@12972.4]
  wire [11:0] _T_617; // @[Cat.scala 30:58:@12974.4]
  wire [11:0] _T_619; // @[Cat.scala 30:58:@12976.4]
  wire [11:0] _T_620; // @[Mux.scala 31:69:@12977.4]
  wire [11:0] _T_621; // @[Mux.scala 31:69:@12978.4]
  wire [11:0] _T_622; // @[Mux.scala 31:69:@12979.4]
  wire [11:0] _T_623; // @[Mux.scala 31:69:@12980.4]
  wire [11:0] _T_624; // @[Mux.scala 31:69:@12981.4]
  wire [11:0] _T_625; // @[Mux.scala 31:69:@12982.4]
  wire [11:0] _T_626; // @[Mux.scala 31:69:@12983.4]
  wire [11:0] _T_627; // @[Mux.scala 31:69:@12984.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@12992.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@12993.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@12996.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@12997.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13000.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13001.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13004.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13005.4]
  wire  _T_658; // @[MemPrimitives.scala 110:210:@13008.4]
  wire  _T_659; // @[MemPrimitives.scala 110:228:@13009.4]
  wire  _T_664; // @[MemPrimitives.scala 110:210:@13012.4]
  wire  _T_665; // @[MemPrimitives.scala 110:228:@13013.4]
  wire  _T_670; // @[MemPrimitives.scala 110:210:@13016.4]
  wire  _T_671; // @[MemPrimitives.scala 110:228:@13017.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@13020.4]
  wire  _T_677; // @[MemPrimitives.scala 110:228:@13021.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13024.4]
  wire  _T_683; // @[MemPrimitives.scala 110:228:@13025.4]
  wire  _T_685; // @[MemPrimitives.scala 126:35:@13039.4]
  wire  _T_686; // @[MemPrimitives.scala 126:35:@13040.4]
  wire  _T_687; // @[MemPrimitives.scala 126:35:@13041.4]
  wire  _T_688; // @[MemPrimitives.scala 126:35:@13042.4]
  wire  _T_689; // @[MemPrimitives.scala 126:35:@13043.4]
  wire  _T_690; // @[MemPrimitives.scala 126:35:@13044.4]
  wire  _T_691; // @[MemPrimitives.scala 126:35:@13045.4]
  wire  _T_692; // @[MemPrimitives.scala 126:35:@13046.4]
  wire  _T_693; // @[MemPrimitives.scala 126:35:@13047.4]
  wire [11:0] _T_695; // @[Cat.scala 30:58:@13049.4]
  wire [11:0] _T_697; // @[Cat.scala 30:58:@13051.4]
  wire [11:0] _T_699; // @[Cat.scala 30:58:@13053.4]
  wire [11:0] _T_701; // @[Cat.scala 30:58:@13055.4]
  wire [11:0] _T_703; // @[Cat.scala 30:58:@13057.4]
  wire [11:0] _T_705; // @[Cat.scala 30:58:@13059.4]
  wire [11:0] _T_707; // @[Cat.scala 30:58:@13061.4]
  wire [11:0] _T_709; // @[Cat.scala 30:58:@13063.4]
  wire [11:0] _T_711; // @[Cat.scala 30:58:@13065.4]
  wire [11:0] _T_712; // @[Mux.scala 31:69:@13066.4]
  wire [11:0] _T_713; // @[Mux.scala 31:69:@13067.4]
  wire [11:0] _T_714; // @[Mux.scala 31:69:@13068.4]
  wire [11:0] _T_715; // @[Mux.scala 31:69:@13069.4]
  wire [11:0] _T_716; // @[Mux.scala 31:69:@13070.4]
  wire [11:0] _T_717; // @[Mux.scala 31:69:@13071.4]
  wire [11:0] _T_718; // @[Mux.scala 31:69:@13072.4]
  wire [11:0] _T_719; // @[Mux.scala 31:69:@13073.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@13080.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@13082.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@13084.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@13086.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@13088.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@13090.4]
  wire  _T_742; // @[MemPrimitives.scala 110:210:@13092.4]
  wire  _T_745; // @[MemPrimitives.scala 110:228:@13094.4]
  wire  _T_748; // @[MemPrimitives.scala 110:210:@13096.4]
  wire  _T_751; // @[MemPrimitives.scala 110:228:@13098.4]
  wire  _T_754; // @[MemPrimitives.scala 110:210:@13100.4]
  wire  _T_757; // @[MemPrimitives.scala 110:228:@13102.4]
  wire  _T_760; // @[MemPrimitives.scala 110:210:@13104.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@13106.4]
  wire  _T_766; // @[MemPrimitives.scala 110:210:@13108.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@13110.4]
  wire  _T_772; // @[MemPrimitives.scala 110:210:@13112.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@13114.4]
  wire  _T_777; // @[MemPrimitives.scala 126:35:@13128.4]
  wire  _T_778; // @[MemPrimitives.scala 126:35:@13129.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@13130.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@13131.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@13132.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@13133.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@13134.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@13135.4]
  wire  _T_785; // @[MemPrimitives.scala 126:35:@13136.4]
  wire [11:0] _T_787; // @[Cat.scala 30:58:@13138.4]
  wire [11:0] _T_789; // @[Cat.scala 30:58:@13140.4]
  wire [11:0] _T_791; // @[Cat.scala 30:58:@13142.4]
  wire [11:0] _T_793; // @[Cat.scala 30:58:@13144.4]
  wire [11:0] _T_795; // @[Cat.scala 30:58:@13146.4]
  wire [11:0] _T_797; // @[Cat.scala 30:58:@13148.4]
  wire [11:0] _T_799; // @[Cat.scala 30:58:@13150.4]
  wire [11:0] _T_801; // @[Cat.scala 30:58:@13152.4]
  wire [11:0] _T_803; // @[Cat.scala 30:58:@13154.4]
  wire [11:0] _T_804; // @[Mux.scala 31:69:@13155.4]
  wire [11:0] _T_805; // @[Mux.scala 31:69:@13156.4]
  wire [11:0] _T_806; // @[Mux.scala 31:69:@13157.4]
  wire [11:0] _T_807; // @[Mux.scala 31:69:@13158.4]
  wire [11:0] _T_808; // @[Mux.scala 31:69:@13159.4]
  wire [11:0] _T_809; // @[Mux.scala 31:69:@13160.4]
  wire [11:0] _T_810; // @[Mux.scala 31:69:@13161.4]
  wire [11:0] _T_811; // @[Mux.scala 31:69:@13162.4]
  wire  _T_819; // @[MemPrimitives.scala 110:228:@13171.4]
  wire  _T_825; // @[MemPrimitives.scala 110:228:@13175.4]
  wire  _T_831; // @[MemPrimitives.scala 110:228:@13179.4]
  wire  _T_837; // @[MemPrimitives.scala 110:228:@13183.4]
  wire  _T_843; // @[MemPrimitives.scala 110:228:@13187.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@13191.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@13195.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@13199.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@13203.4]
  wire  _T_869; // @[MemPrimitives.scala 126:35:@13217.4]
  wire  _T_870; // @[MemPrimitives.scala 126:35:@13218.4]
  wire  _T_871; // @[MemPrimitives.scala 126:35:@13219.4]
  wire  _T_872; // @[MemPrimitives.scala 126:35:@13220.4]
  wire  _T_873; // @[MemPrimitives.scala 126:35:@13221.4]
  wire  _T_874; // @[MemPrimitives.scala 126:35:@13222.4]
  wire  _T_875; // @[MemPrimitives.scala 126:35:@13223.4]
  wire  _T_876; // @[MemPrimitives.scala 126:35:@13224.4]
  wire  _T_877; // @[MemPrimitives.scala 126:35:@13225.4]
  wire [11:0] _T_879; // @[Cat.scala 30:58:@13227.4]
  wire [11:0] _T_881; // @[Cat.scala 30:58:@13229.4]
  wire [11:0] _T_883; // @[Cat.scala 30:58:@13231.4]
  wire [11:0] _T_885; // @[Cat.scala 30:58:@13233.4]
  wire [11:0] _T_887; // @[Cat.scala 30:58:@13235.4]
  wire [11:0] _T_889; // @[Cat.scala 30:58:@13237.4]
  wire [11:0] _T_891; // @[Cat.scala 30:58:@13239.4]
  wire [11:0] _T_893; // @[Cat.scala 30:58:@13241.4]
  wire [11:0] _T_895; // @[Cat.scala 30:58:@13243.4]
  wire [11:0] _T_896; // @[Mux.scala 31:69:@13244.4]
  wire [11:0] _T_897; // @[Mux.scala 31:69:@13245.4]
  wire [11:0] _T_898; // @[Mux.scala 31:69:@13246.4]
  wire [11:0] _T_899; // @[Mux.scala 31:69:@13247.4]
  wire [11:0] _T_900; // @[Mux.scala 31:69:@13248.4]
  wire [11:0] _T_901; // @[Mux.scala 31:69:@13249.4]
  wire [11:0] _T_902; // @[Mux.scala 31:69:@13250.4]
  wire [11:0] _T_903; // @[Mux.scala 31:69:@13251.4]
  wire  _T_911; // @[MemPrimitives.scala 110:228:@13260.4]
  wire  _T_917; // @[MemPrimitives.scala 110:228:@13264.4]
  wire  _T_923; // @[MemPrimitives.scala 110:228:@13268.4]
  wire  _T_929; // @[MemPrimitives.scala 110:228:@13272.4]
  wire  _T_935; // @[MemPrimitives.scala 110:228:@13276.4]
  wire  _T_941; // @[MemPrimitives.scala 110:228:@13280.4]
  wire  _T_947; // @[MemPrimitives.scala 110:228:@13284.4]
  wire  _T_953; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_959; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_961; // @[MemPrimitives.scala 126:35:@13306.4]
  wire  _T_962; // @[MemPrimitives.scala 126:35:@13307.4]
  wire  _T_963; // @[MemPrimitives.scala 126:35:@13308.4]
  wire  _T_964; // @[MemPrimitives.scala 126:35:@13309.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13310.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13311.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13312.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13313.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13314.4]
  wire [11:0] _T_971; // @[Cat.scala 30:58:@13316.4]
  wire [11:0] _T_973; // @[Cat.scala 30:58:@13318.4]
  wire [11:0] _T_975; // @[Cat.scala 30:58:@13320.4]
  wire [11:0] _T_977; // @[Cat.scala 30:58:@13322.4]
  wire [11:0] _T_979; // @[Cat.scala 30:58:@13324.4]
  wire [11:0] _T_981; // @[Cat.scala 30:58:@13326.4]
  wire [11:0] _T_983; // @[Cat.scala 30:58:@13328.4]
  wire [11:0] _T_985; // @[Cat.scala 30:58:@13330.4]
  wire [11:0] _T_987; // @[Cat.scala 30:58:@13332.4]
  wire [11:0] _T_988; // @[Mux.scala 31:69:@13333.4]
  wire [11:0] _T_989; // @[Mux.scala 31:69:@13334.4]
  wire [11:0] _T_990; // @[Mux.scala 31:69:@13335.4]
  wire [11:0] _T_991; // @[Mux.scala 31:69:@13336.4]
  wire [11:0] _T_992; // @[Mux.scala 31:69:@13337.4]
  wire [11:0] _T_993; // @[Mux.scala 31:69:@13338.4]
  wire [11:0] _T_994; // @[Mux.scala 31:69:@13339.4]
  wire [11:0] _T_995; // @[Mux.scala 31:69:@13340.4]
  wire  _T_1000; // @[MemPrimitives.scala 110:210:@13347.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@13349.4]
  wire  _T_1006; // @[MemPrimitives.scala 110:210:@13351.4]
  wire  _T_1009; // @[MemPrimitives.scala 110:228:@13353.4]
  wire  _T_1012; // @[MemPrimitives.scala 110:210:@13355.4]
  wire  _T_1015; // @[MemPrimitives.scala 110:228:@13357.4]
  wire  _T_1018; // @[MemPrimitives.scala 110:210:@13359.4]
  wire  _T_1021; // @[MemPrimitives.scala 110:228:@13361.4]
  wire  _T_1024; // @[MemPrimitives.scala 110:210:@13363.4]
  wire  _T_1027; // @[MemPrimitives.scala 110:228:@13365.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@13367.4]
  wire  _T_1033; // @[MemPrimitives.scala 110:228:@13369.4]
  wire  _T_1036; // @[MemPrimitives.scala 110:210:@13371.4]
  wire  _T_1039; // @[MemPrimitives.scala 110:228:@13373.4]
  wire  _T_1042; // @[MemPrimitives.scala 110:210:@13375.4]
  wire  _T_1045; // @[MemPrimitives.scala 110:228:@13377.4]
  wire  _T_1048; // @[MemPrimitives.scala 110:210:@13379.4]
  wire  _T_1051; // @[MemPrimitives.scala 110:228:@13381.4]
  wire  _T_1053; // @[MemPrimitives.scala 126:35:@13395.4]
  wire  _T_1054; // @[MemPrimitives.scala 126:35:@13396.4]
  wire  _T_1055; // @[MemPrimitives.scala 126:35:@13397.4]
  wire  _T_1056; // @[MemPrimitives.scala 126:35:@13398.4]
  wire  _T_1057; // @[MemPrimitives.scala 126:35:@13399.4]
  wire  _T_1058; // @[MemPrimitives.scala 126:35:@13400.4]
  wire  _T_1059; // @[MemPrimitives.scala 126:35:@13401.4]
  wire  _T_1060; // @[MemPrimitives.scala 126:35:@13402.4]
  wire  _T_1061; // @[MemPrimitives.scala 126:35:@13403.4]
  wire [11:0] _T_1063; // @[Cat.scala 30:58:@13405.4]
  wire [11:0] _T_1065; // @[Cat.scala 30:58:@13407.4]
  wire [11:0] _T_1067; // @[Cat.scala 30:58:@13409.4]
  wire [11:0] _T_1069; // @[Cat.scala 30:58:@13411.4]
  wire [11:0] _T_1071; // @[Cat.scala 30:58:@13413.4]
  wire [11:0] _T_1073; // @[Cat.scala 30:58:@13415.4]
  wire [11:0] _T_1075; // @[Cat.scala 30:58:@13417.4]
  wire [11:0] _T_1077; // @[Cat.scala 30:58:@13419.4]
  wire [11:0] _T_1079; // @[Cat.scala 30:58:@13421.4]
  wire [11:0] _T_1080; // @[Mux.scala 31:69:@13422.4]
  wire [11:0] _T_1081; // @[Mux.scala 31:69:@13423.4]
  wire [11:0] _T_1082; // @[Mux.scala 31:69:@13424.4]
  wire [11:0] _T_1083; // @[Mux.scala 31:69:@13425.4]
  wire [11:0] _T_1084; // @[Mux.scala 31:69:@13426.4]
  wire [11:0] _T_1085; // @[Mux.scala 31:69:@13427.4]
  wire [11:0] _T_1086; // @[Mux.scala 31:69:@13428.4]
  wire [11:0] _T_1087; // @[Mux.scala 31:69:@13429.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@13438.4]
  wire  _T_1101; // @[MemPrimitives.scala 110:228:@13442.4]
  wire  _T_1107; // @[MemPrimitives.scala 110:228:@13446.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:228:@13450.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13454.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13458.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13462.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13466.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13470.4]
  wire  _T_1145; // @[MemPrimitives.scala 126:35:@13484.4]
  wire  _T_1146; // @[MemPrimitives.scala 126:35:@13485.4]
  wire  _T_1147; // @[MemPrimitives.scala 126:35:@13486.4]
  wire  _T_1148; // @[MemPrimitives.scala 126:35:@13487.4]
  wire  _T_1149; // @[MemPrimitives.scala 126:35:@13488.4]
  wire  _T_1150; // @[MemPrimitives.scala 126:35:@13489.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13490.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13491.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13492.4]
  wire [11:0] _T_1155; // @[Cat.scala 30:58:@13494.4]
  wire [11:0] _T_1157; // @[Cat.scala 30:58:@13496.4]
  wire [11:0] _T_1159; // @[Cat.scala 30:58:@13498.4]
  wire [11:0] _T_1161; // @[Cat.scala 30:58:@13500.4]
  wire [11:0] _T_1163; // @[Cat.scala 30:58:@13502.4]
  wire [11:0] _T_1165; // @[Cat.scala 30:58:@13504.4]
  wire [11:0] _T_1167; // @[Cat.scala 30:58:@13506.4]
  wire [11:0] _T_1169; // @[Cat.scala 30:58:@13508.4]
  wire [11:0] _T_1171; // @[Cat.scala 30:58:@13510.4]
  wire [11:0] _T_1172; // @[Mux.scala 31:69:@13511.4]
  wire [11:0] _T_1173; // @[Mux.scala 31:69:@13512.4]
  wire [11:0] _T_1174; // @[Mux.scala 31:69:@13513.4]
  wire [11:0] _T_1175; // @[Mux.scala 31:69:@13514.4]
  wire [11:0] _T_1176; // @[Mux.scala 31:69:@13515.4]
  wire [11:0] _T_1177; // @[Mux.scala 31:69:@13516.4]
  wire [11:0] _T_1178; // @[Mux.scala 31:69:@13517.4]
  wire [11:0] _T_1179; // @[Mux.scala 31:69:@13518.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13527.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13531.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13535.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13539.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13543.4]
  wire  _T_1217; // @[MemPrimitives.scala 110:228:@13547.4]
  wire  _T_1223; // @[MemPrimitives.scala 110:228:@13551.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:228:@13555.4]
  wire  _T_1235; // @[MemPrimitives.scala 110:228:@13559.4]
  wire  _T_1237; // @[MemPrimitives.scala 126:35:@13573.4]
  wire  _T_1238; // @[MemPrimitives.scala 126:35:@13574.4]
  wire  _T_1239; // @[MemPrimitives.scala 126:35:@13575.4]
  wire  _T_1240; // @[MemPrimitives.scala 126:35:@13576.4]
  wire  _T_1241; // @[MemPrimitives.scala 126:35:@13577.4]
  wire  _T_1242; // @[MemPrimitives.scala 126:35:@13578.4]
  wire  _T_1243; // @[MemPrimitives.scala 126:35:@13579.4]
  wire  _T_1244; // @[MemPrimitives.scala 126:35:@13580.4]
  wire  _T_1245; // @[MemPrimitives.scala 126:35:@13581.4]
  wire [11:0] _T_1247; // @[Cat.scala 30:58:@13583.4]
  wire [11:0] _T_1249; // @[Cat.scala 30:58:@13585.4]
  wire [11:0] _T_1251; // @[Cat.scala 30:58:@13587.4]
  wire [11:0] _T_1253; // @[Cat.scala 30:58:@13589.4]
  wire [11:0] _T_1255; // @[Cat.scala 30:58:@13591.4]
  wire [11:0] _T_1257; // @[Cat.scala 30:58:@13593.4]
  wire [11:0] _T_1259; // @[Cat.scala 30:58:@13595.4]
  wire [11:0] _T_1261; // @[Cat.scala 30:58:@13597.4]
  wire [11:0] _T_1263; // @[Cat.scala 30:58:@13599.4]
  wire [11:0] _T_1264; // @[Mux.scala 31:69:@13600.4]
  wire [11:0] _T_1265; // @[Mux.scala 31:69:@13601.4]
  wire [11:0] _T_1266; // @[Mux.scala 31:69:@13602.4]
  wire [11:0] _T_1267; // @[Mux.scala 31:69:@13603.4]
  wire [11:0] _T_1268; // @[Mux.scala 31:69:@13604.4]
  wire [11:0] _T_1269; // @[Mux.scala 31:69:@13605.4]
  wire [11:0] _T_1270; // @[Mux.scala 31:69:@13606.4]
  wire [11:0] _T_1271; // @[Mux.scala 31:69:@13607.4]
  wire  _T_1276; // @[MemPrimitives.scala 110:210:@13614.4]
  wire  _T_1279; // @[MemPrimitives.scala 110:228:@13616.4]
  wire  _T_1282; // @[MemPrimitives.scala 110:210:@13618.4]
  wire  _T_1285; // @[MemPrimitives.scala 110:228:@13620.4]
  wire  _T_1288; // @[MemPrimitives.scala 110:210:@13622.4]
  wire  _T_1291; // @[MemPrimitives.scala 110:228:@13624.4]
  wire  _T_1294; // @[MemPrimitives.scala 110:210:@13626.4]
  wire  _T_1297; // @[MemPrimitives.scala 110:228:@13628.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@13630.4]
  wire  _T_1303; // @[MemPrimitives.scala 110:228:@13632.4]
  wire  _T_1306; // @[MemPrimitives.scala 110:210:@13634.4]
  wire  _T_1309; // @[MemPrimitives.scala 110:228:@13636.4]
  wire  _T_1312; // @[MemPrimitives.scala 110:210:@13638.4]
  wire  _T_1315; // @[MemPrimitives.scala 110:228:@13640.4]
  wire  _T_1318; // @[MemPrimitives.scala 110:210:@13642.4]
  wire  _T_1321; // @[MemPrimitives.scala 110:228:@13644.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@13646.4]
  wire  _T_1327; // @[MemPrimitives.scala 110:228:@13648.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@13662.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@13663.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@13664.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@13665.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@13666.4]
  wire  _T_1334; // @[MemPrimitives.scala 126:35:@13667.4]
  wire  _T_1335; // @[MemPrimitives.scala 126:35:@13668.4]
  wire  _T_1336; // @[MemPrimitives.scala 126:35:@13669.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13670.4]
  wire [11:0] _T_1339; // @[Cat.scala 30:58:@13672.4]
  wire [11:0] _T_1341; // @[Cat.scala 30:58:@13674.4]
  wire [11:0] _T_1343; // @[Cat.scala 30:58:@13676.4]
  wire [11:0] _T_1345; // @[Cat.scala 30:58:@13678.4]
  wire [11:0] _T_1347; // @[Cat.scala 30:58:@13680.4]
  wire [11:0] _T_1349; // @[Cat.scala 30:58:@13682.4]
  wire [11:0] _T_1351; // @[Cat.scala 30:58:@13684.4]
  wire [11:0] _T_1353; // @[Cat.scala 30:58:@13686.4]
  wire [11:0] _T_1355; // @[Cat.scala 30:58:@13688.4]
  wire [11:0] _T_1356; // @[Mux.scala 31:69:@13689.4]
  wire [11:0] _T_1357; // @[Mux.scala 31:69:@13690.4]
  wire [11:0] _T_1358; // @[Mux.scala 31:69:@13691.4]
  wire [11:0] _T_1359; // @[Mux.scala 31:69:@13692.4]
  wire [11:0] _T_1360; // @[Mux.scala 31:69:@13693.4]
  wire [11:0] _T_1361; // @[Mux.scala 31:69:@13694.4]
  wire [11:0] _T_1362; // @[Mux.scala 31:69:@13695.4]
  wire [11:0] _T_1363; // @[Mux.scala 31:69:@13696.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@13705.4]
  wire  _T_1377; // @[MemPrimitives.scala 110:228:@13709.4]
  wire  _T_1383; // @[MemPrimitives.scala 110:228:@13713.4]
  wire  _T_1389; // @[MemPrimitives.scala 110:228:@13717.4]
  wire  _T_1395; // @[MemPrimitives.scala 110:228:@13721.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:228:@13725.4]
  wire  _T_1407; // @[MemPrimitives.scala 110:228:@13729.4]
  wire  _T_1413; // @[MemPrimitives.scala 110:228:@13733.4]
  wire  _T_1419; // @[MemPrimitives.scala 110:228:@13737.4]
  wire  _T_1421; // @[MemPrimitives.scala 126:35:@13751.4]
  wire  _T_1422; // @[MemPrimitives.scala 126:35:@13752.4]
  wire  _T_1423; // @[MemPrimitives.scala 126:35:@13753.4]
  wire  _T_1424; // @[MemPrimitives.scala 126:35:@13754.4]
  wire  _T_1425; // @[MemPrimitives.scala 126:35:@13755.4]
  wire  _T_1426; // @[MemPrimitives.scala 126:35:@13756.4]
  wire  _T_1427; // @[MemPrimitives.scala 126:35:@13757.4]
  wire  _T_1428; // @[MemPrimitives.scala 126:35:@13758.4]
  wire  _T_1429; // @[MemPrimitives.scala 126:35:@13759.4]
  wire [11:0] _T_1431; // @[Cat.scala 30:58:@13761.4]
  wire [11:0] _T_1433; // @[Cat.scala 30:58:@13763.4]
  wire [11:0] _T_1435; // @[Cat.scala 30:58:@13765.4]
  wire [11:0] _T_1437; // @[Cat.scala 30:58:@13767.4]
  wire [11:0] _T_1439; // @[Cat.scala 30:58:@13769.4]
  wire [11:0] _T_1441; // @[Cat.scala 30:58:@13771.4]
  wire [11:0] _T_1443; // @[Cat.scala 30:58:@13773.4]
  wire [11:0] _T_1445; // @[Cat.scala 30:58:@13775.4]
  wire [11:0] _T_1447; // @[Cat.scala 30:58:@13777.4]
  wire [11:0] _T_1448; // @[Mux.scala 31:69:@13778.4]
  wire [11:0] _T_1449; // @[Mux.scala 31:69:@13779.4]
  wire [11:0] _T_1450; // @[Mux.scala 31:69:@13780.4]
  wire [11:0] _T_1451; // @[Mux.scala 31:69:@13781.4]
  wire [11:0] _T_1452; // @[Mux.scala 31:69:@13782.4]
  wire [11:0] _T_1453; // @[Mux.scala 31:69:@13783.4]
  wire [11:0] _T_1454; // @[Mux.scala 31:69:@13784.4]
  wire [11:0] _T_1455; // @[Mux.scala 31:69:@13785.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@13794.4]
  wire  _T_1469; // @[MemPrimitives.scala 110:228:@13798.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:228:@13802.4]
  wire  _T_1481; // @[MemPrimitives.scala 110:228:@13806.4]
  wire  _T_1487; // @[MemPrimitives.scala 110:228:@13810.4]
  wire  _T_1493; // @[MemPrimitives.scala 110:228:@13814.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:228:@13818.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:228:@13822.4]
  wire  _T_1511; // @[MemPrimitives.scala 110:228:@13826.4]
  wire  _T_1513; // @[MemPrimitives.scala 126:35:@13840.4]
  wire  _T_1514; // @[MemPrimitives.scala 126:35:@13841.4]
  wire  _T_1515; // @[MemPrimitives.scala 126:35:@13842.4]
  wire  _T_1516; // @[MemPrimitives.scala 126:35:@13843.4]
  wire  _T_1517; // @[MemPrimitives.scala 126:35:@13844.4]
  wire  _T_1518; // @[MemPrimitives.scala 126:35:@13845.4]
  wire  _T_1519; // @[MemPrimitives.scala 126:35:@13846.4]
  wire  _T_1520; // @[MemPrimitives.scala 126:35:@13847.4]
  wire  _T_1521; // @[MemPrimitives.scala 126:35:@13848.4]
  wire [11:0] _T_1523; // @[Cat.scala 30:58:@13850.4]
  wire [11:0] _T_1525; // @[Cat.scala 30:58:@13852.4]
  wire [11:0] _T_1527; // @[Cat.scala 30:58:@13854.4]
  wire [11:0] _T_1529; // @[Cat.scala 30:58:@13856.4]
  wire [11:0] _T_1531; // @[Cat.scala 30:58:@13858.4]
  wire [11:0] _T_1533; // @[Cat.scala 30:58:@13860.4]
  wire [11:0] _T_1535; // @[Cat.scala 30:58:@13862.4]
  wire [11:0] _T_1537; // @[Cat.scala 30:58:@13864.4]
  wire [11:0] _T_1539; // @[Cat.scala 30:58:@13866.4]
  wire [11:0] _T_1540; // @[Mux.scala 31:69:@13867.4]
  wire [11:0] _T_1541; // @[Mux.scala 31:69:@13868.4]
  wire [11:0] _T_1542; // @[Mux.scala 31:69:@13869.4]
  wire [11:0] _T_1543; // @[Mux.scala 31:69:@13870.4]
  wire [11:0] _T_1544; // @[Mux.scala 31:69:@13871.4]
  wire [11:0] _T_1545; // @[Mux.scala 31:69:@13872.4]
  wire [11:0] _T_1546; // @[Mux.scala 31:69:@13873.4]
  wire [11:0] _T_1547; // @[Mux.scala 31:69:@13874.4]
  wire  _T_1643; // @[package.scala 96:25:@14003.4 package.scala 96:25:@14004.4]
  wire [31:0] _T_1647; // @[Mux.scala 31:69:@14013.4]
  wire  _T_1640; // @[package.scala 96:25:@13995.4 package.scala 96:25:@13996.4]
  wire [31:0] _T_1648; // @[Mux.scala 31:69:@14014.4]
  wire  _T_1637; // @[package.scala 96:25:@13987.4 package.scala 96:25:@13988.4]
  wire [31:0] _T_1649; // @[Mux.scala 31:69:@14015.4]
  wire  _T_1634; // @[package.scala 96:25:@13979.4 package.scala 96:25:@13980.4]
  wire [31:0] _T_1650; // @[Mux.scala 31:69:@14016.4]
  wire  _T_1631; // @[package.scala 96:25:@13971.4 package.scala 96:25:@13972.4]
  wire [31:0] _T_1651; // @[Mux.scala 31:69:@14017.4]
  wire  _T_1628; // @[package.scala 96:25:@13963.4 package.scala 96:25:@13964.4]
  wire [31:0] _T_1652; // @[Mux.scala 31:69:@14018.4]
  wire  _T_1625; // @[package.scala 96:25:@13955.4 package.scala 96:25:@13956.4]
  wire [31:0] _T_1653; // @[Mux.scala 31:69:@14019.4]
  wire  _T_1622; // @[package.scala 96:25:@13947.4 package.scala 96:25:@13948.4]
  wire [31:0] _T_1654; // @[Mux.scala 31:69:@14020.4]
  wire  _T_1619; // @[package.scala 96:25:@13939.4 package.scala 96:25:@13940.4]
  wire [31:0] _T_1655; // @[Mux.scala 31:69:@14021.4]
  wire  _T_1616; // @[package.scala 96:25:@13931.4 package.scala 96:25:@13932.4]
  wire [31:0] _T_1656; // @[Mux.scala 31:69:@14022.4]
  wire  _T_1613; // @[package.scala 96:25:@13923.4 package.scala 96:25:@13924.4]
  wire  _T_1750; // @[package.scala 96:25:@14147.4 package.scala 96:25:@14148.4]
  wire [31:0] _T_1754; // @[Mux.scala 31:69:@14157.4]
  wire  _T_1747; // @[package.scala 96:25:@14139.4 package.scala 96:25:@14140.4]
  wire [31:0] _T_1755; // @[Mux.scala 31:69:@14158.4]
  wire  _T_1744; // @[package.scala 96:25:@14131.4 package.scala 96:25:@14132.4]
  wire [31:0] _T_1756; // @[Mux.scala 31:69:@14159.4]
  wire  _T_1741; // @[package.scala 96:25:@14123.4 package.scala 96:25:@14124.4]
  wire [31:0] _T_1757; // @[Mux.scala 31:69:@14160.4]
  wire  _T_1738; // @[package.scala 96:25:@14115.4 package.scala 96:25:@14116.4]
  wire [31:0] _T_1758; // @[Mux.scala 31:69:@14161.4]
  wire  _T_1735; // @[package.scala 96:25:@14107.4 package.scala 96:25:@14108.4]
  wire [31:0] _T_1759; // @[Mux.scala 31:69:@14162.4]
  wire  _T_1732; // @[package.scala 96:25:@14099.4 package.scala 96:25:@14100.4]
  wire [31:0] _T_1760; // @[Mux.scala 31:69:@14163.4]
  wire  _T_1729; // @[package.scala 96:25:@14091.4 package.scala 96:25:@14092.4]
  wire [31:0] _T_1761; // @[Mux.scala 31:69:@14164.4]
  wire  _T_1726; // @[package.scala 96:25:@14083.4 package.scala 96:25:@14084.4]
  wire [31:0] _T_1762; // @[Mux.scala 31:69:@14165.4]
  wire  _T_1723; // @[package.scala 96:25:@14075.4 package.scala 96:25:@14076.4]
  wire [31:0] _T_1763; // @[Mux.scala 31:69:@14166.4]
  wire  _T_1720; // @[package.scala 96:25:@14067.4 package.scala 96:25:@14068.4]
  wire  _T_1857; // @[package.scala 96:25:@14291.4 package.scala 96:25:@14292.4]
  wire [31:0] _T_1861; // @[Mux.scala 31:69:@14301.4]
  wire  _T_1854; // @[package.scala 96:25:@14283.4 package.scala 96:25:@14284.4]
  wire [31:0] _T_1862; // @[Mux.scala 31:69:@14302.4]
  wire  _T_1851; // @[package.scala 96:25:@14275.4 package.scala 96:25:@14276.4]
  wire [31:0] _T_1863; // @[Mux.scala 31:69:@14303.4]
  wire  _T_1848; // @[package.scala 96:25:@14267.4 package.scala 96:25:@14268.4]
  wire [31:0] _T_1864; // @[Mux.scala 31:69:@14304.4]
  wire  _T_1845; // @[package.scala 96:25:@14259.4 package.scala 96:25:@14260.4]
  wire [31:0] _T_1865; // @[Mux.scala 31:69:@14305.4]
  wire  _T_1842; // @[package.scala 96:25:@14251.4 package.scala 96:25:@14252.4]
  wire [31:0] _T_1866; // @[Mux.scala 31:69:@14306.4]
  wire  _T_1839; // @[package.scala 96:25:@14243.4 package.scala 96:25:@14244.4]
  wire [31:0] _T_1867; // @[Mux.scala 31:69:@14307.4]
  wire  _T_1836; // @[package.scala 96:25:@14235.4 package.scala 96:25:@14236.4]
  wire [31:0] _T_1868; // @[Mux.scala 31:69:@14308.4]
  wire  _T_1833; // @[package.scala 96:25:@14227.4 package.scala 96:25:@14228.4]
  wire [31:0] _T_1869; // @[Mux.scala 31:69:@14309.4]
  wire  _T_1830; // @[package.scala 96:25:@14219.4 package.scala 96:25:@14220.4]
  wire [31:0] _T_1870; // @[Mux.scala 31:69:@14310.4]
  wire  _T_1827; // @[package.scala 96:25:@14211.4 package.scala 96:25:@14212.4]
  wire  _T_1964; // @[package.scala 96:25:@14435.4 package.scala 96:25:@14436.4]
  wire [31:0] _T_1968; // @[Mux.scala 31:69:@14445.4]
  wire  _T_1961; // @[package.scala 96:25:@14427.4 package.scala 96:25:@14428.4]
  wire [31:0] _T_1969; // @[Mux.scala 31:69:@14446.4]
  wire  _T_1958; // @[package.scala 96:25:@14419.4 package.scala 96:25:@14420.4]
  wire [31:0] _T_1970; // @[Mux.scala 31:69:@14447.4]
  wire  _T_1955; // @[package.scala 96:25:@14411.4 package.scala 96:25:@14412.4]
  wire [31:0] _T_1971; // @[Mux.scala 31:69:@14448.4]
  wire  _T_1952; // @[package.scala 96:25:@14403.4 package.scala 96:25:@14404.4]
  wire [31:0] _T_1972; // @[Mux.scala 31:69:@14449.4]
  wire  _T_1949; // @[package.scala 96:25:@14395.4 package.scala 96:25:@14396.4]
  wire [31:0] _T_1973; // @[Mux.scala 31:69:@14450.4]
  wire  _T_1946; // @[package.scala 96:25:@14387.4 package.scala 96:25:@14388.4]
  wire [31:0] _T_1974; // @[Mux.scala 31:69:@14451.4]
  wire  _T_1943; // @[package.scala 96:25:@14379.4 package.scala 96:25:@14380.4]
  wire [31:0] _T_1975; // @[Mux.scala 31:69:@14452.4]
  wire  _T_1940; // @[package.scala 96:25:@14371.4 package.scala 96:25:@14372.4]
  wire [31:0] _T_1976; // @[Mux.scala 31:69:@14453.4]
  wire  _T_1937; // @[package.scala 96:25:@14363.4 package.scala 96:25:@14364.4]
  wire [31:0] _T_1977; // @[Mux.scala 31:69:@14454.4]
  wire  _T_1934; // @[package.scala 96:25:@14355.4 package.scala 96:25:@14356.4]
  wire  _T_2071; // @[package.scala 96:25:@14579.4 package.scala 96:25:@14580.4]
  wire [31:0] _T_2075; // @[Mux.scala 31:69:@14589.4]
  wire  _T_2068; // @[package.scala 96:25:@14571.4 package.scala 96:25:@14572.4]
  wire [31:0] _T_2076; // @[Mux.scala 31:69:@14590.4]
  wire  _T_2065; // @[package.scala 96:25:@14563.4 package.scala 96:25:@14564.4]
  wire [31:0] _T_2077; // @[Mux.scala 31:69:@14591.4]
  wire  _T_2062; // @[package.scala 96:25:@14555.4 package.scala 96:25:@14556.4]
  wire [31:0] _T_2078; // @[Mux.scala 31:69:@14592.4]
  wire  _T_2059; // @[package.scala 96:25:@14547.4 package.scala 96:25:@14548.4]
  wire [31:0] _T_2079; // @[Mux.scala 31:69:@14593.4]
  wire  _T_2056; // @[package.scala 96:25:@14539.4 package.scala 96:25:@14540.4]
  wire [31:0] _T_2080; // @[Mux.scala 31:69:@14594.4]
  wire  _T_2053; // @[package.scala 96:25:@14531.4 package.scala 96:25:@14532.4]
  wire [31:0] _T_2081; // @[Mux.scala 31:69:@14595.4]
  wire  _T_2050; // @[package.scala 96:25:@14523.4 package.scala 96:25:@14524.4]
  wire [31:0] _T_2082; // @[Mux.scala 31:69:@14596.4]
  wire  _T_2047; // @[package.scala 96:25:@14515.4 package.scala 96:25:@14516.4]
  wire [31:0] _T_2083; // @[Mux.scala 31:69:@14597.4]
  wire  _T_2044; // @[package.scala 96:25:@14507.4 package.scala 96:25:@14508.4]
  wire [31:0] _T_2084; // @[Mux.scala 31:69:@14598.4]
  wire  _T_2041; // @[package.scala 96:25:@14499.4 package.scala 96:25:@14500.4]
  wire  _T_2178; // @[package.scala 96:25:@14723.4 package.scala 96:25:@14724.4]
  wire [31:0] _T_2182; // @[Mux.scala 31:69:@14733.4]
  wire  _T_2175; // @[package.scala 96:25:@14715.4 package.scala 96:25:@14716.4]
  wire [31:0] _T_2183; // @[Mux.scala 31:69:@14734.4]
  wire  _T_2172; // @[package.scala 96:25:@14707.4 package.scala 96:25:@14708.4]
  wire [31:0] _T_2184; // @[Mux.scala 31:69:@14735.4]
  wire  _T_2169; // @[package.scala 96:25:@14699.4 package.scala 96:25:@14700.4]
  wire [31:0] _T_2185; // @[Mux.scala 31:69:@14736.4]
  wire  _T_2166; // @[package.scala 96:25:@14691.4 package.scala 96:25:@14692.4]
  wire [31:0] _T_2186; // @[Mux.scala 31:69:@14737.4]
  wire  _T_2163; // @[package.scala 96:25:@14683.4 package.scala 96:25:@14684.4]
  wire [31:0] _T_2187; // @[Mux.scala 31:69:@14738.4]
  wire  _T_2160; // @[package.scala 96:25:@14675.4 package.scala 96:25:@14676.4]
  wire [31:0] _T_2188; // @[Mux.scala 31:69:@14739.4]
  wire  _T_2157; // @[package.scala 96:25:@14667.4 package.scala 96:25:@14668.4]
  wire [31:0] _T_2189; // @[Mux.scala 31:69:@14740.4]
  wire  _T_2154; // @[package.scala 96:25:@14659.4 package.scala 96:25:@14660.4]
  wire [31:0] _T_2190; // @[Mux.scala 31:69:@14741.4]
  wire  _T_2151; // @[package.scala 96:25:@14651.4 package.scala 96:25:@14652.4]
  wire [31:0] _T_2191; // @[Mux.scala 31:69:@14742.4]
  wire  _T_2148; // @[package.scala 96:25:@14643.4 package.scala 96:25:@14644.4]
  wire  _T_2285; // @[package.scala 96:25:@14867.4 package.scala 96:25:@14868.4]
  wire [31:0] _T_2289; // @[Mux.scala 31:69:@14877.4]
  wire  _T_2282; // @[package.scala 96:25:@14859.4 package.scala 96:25:@14860.4]
  wire [31:0] _T_2290; // @[Mux.scala 31:69:@14878.4]
  wire  _T_2279; // @[package.scala 96:25:@14851.4 package.scala 96:25:@14852.4]
  wire [31:0] _T_2291; // @[Mux.scala 31:69:@14879.4]
  wire  _T_2276; // @[package.scala 96:25:@14843.4 package.scala 96:25:@14844.4]
  wire [31:0] _T_2292; // @[Mux.scala 31:69:@14880.4]
  wire  _T_2273; // @[package.scala 96:25:@14835.4 package.scala 96:25:@14836.4]
  wire [31:0] _T_2293; // @[Mux.scala 31:69:@14881.4]
  wire  _T_2270; // @[package.scala 96:25:@14827.4 package.scala 96:25:@14828.4]
  wire [31:0] _T_2294; // @[Mux.scala 31:69:@14882.4]
  wire  _T_2267; // @[package.scala 96:25:@14819.4 package.scala 96:25:@14820.4]
  wire [31:0] _T_2295; // @[Mux.scala 31:69:@14883.4]
  wire  _T_2264; // @[package.scala 96:25:@14811.4 package.scala 96:25:@14812.4]
  wire [31:0] _T_2296; // @[Mux.scala 31:69:@14884.4]
  wire  _T_2261; // @[package.scala 96:25:@14803.4 package.scala 96:25:@14804.4]
  wire [31:0] _T_2297; // @[Mux.scala 31:69:@14885.4]
  wire  _T_2258; // @[package.scala 96:25:@14795.4 package.scala 96:25:@14796.4]
  wire [31:0] _T_2298; // @[Mux.scala 31:69:@14886.4]
  wire  _T_2255; // @[package.scala 96:25:@14787.4 package.scala 96:25:@14788.4]
  wire  _T_2392; // @[package.scala 96:25:@15011.4 package.scala 96:25:@15012.4]
  wire [31:0] _T_2396; // @[Mux.scala 31:69:@15021.4]
  wire  _T_2389; // @[package.scala 96:25:@15003.4 package.scala 96:25:@15004.4]
  wire [31:0] _T_2397; // @[Mux.scala 31:69:@15022.4]
  wire  _T_2386; // @[package.scala 96:25:@14995.4 package.scala 96:25:@14996.4]
  wire [31:0] _T_2398; // @[Mux.scala 31:69:@15023.4]
  wire  _T_2383; // @[package.scala 96:25:@14987.4 package.scala 96:25:@14988.4]
  wire [31:0] _T_2399; // @[Mux.scala 31:69:@15024.4]
  wire  _T_2380; // @[package.scala 96:25:@14979.4 package.scala 96:25:@14980.4]
  wire [31:0] _T_2400; // @[Mux.scala 31:69:@15025.4]
  wire  _T_2377; // @[package.scala 96:25:@14971.4 package.scala 96:25:@14972.4]
  wire [31:0] _T_2401; // @[Mux.scala 31:69:@15026.4]
  wire  _T_2374; // @[package.scala 96:25:@14963.4 package.scala 96:25:@14964.4]
  wire [31:0] _T_2402; // @[Mux.scala 31:69:@15027.4]
  wire  _T_2371; // @[package.scala 96:25:@14955.4 package.scala 96:25:@14956.4]
  wire [31:0] _T_2403; // @[Mux.scala 31:69:@15028.4]
  wire  _T_2368; // @[package.scala 96:25:@14947.4 package.scala 96:25:@14948.4]
  wire [31:0] _T_2404; // @[Mux.scala 31:69:@15029.4]
  wire  _T_2365; // @[package.scala 96:25:@14939.4 package.scala 96:25:@14940.4]
  wire [31:0] _T_2405; // @[Mux.scala 31:69:@15030.4]
  wire  _T_2362; // @[package.scala 96:25:@14931.4 package.scala 96:25:@14932.4]
  wire  _T_2499; // @[package.scala 96:25:@15155.4 package.scala 96:25:@15156.4]
  wire [31:0] _T_2503; // @[Mux.scala 31:69:@15165.4]
  wire  _T_2496; // @[package.scala 96:25:@15147.4 package.scala 96:25:@15148.4]
  wire [31:0] _T_2504; // @[Mux.scala 31:69:@15166.4]
  wire  _T_2493; // @[package.scala 96:25:@15139.4 package.scala 96:25:@15140.4]
  wire [31:0] _T_2505; // @[Mux.scala 31:69:@15167.4]
  wire  _T_2490; // @[package.scala 96:25:@15131.4 package.scala 96:25:@15132.4]
  wire [31:0] _T_2506; // @[Mux.scala 31:69:@15168.4]
  wire  _T_2487; // @[package.scala 96:25:@15123.4 package.scala 96:25:@15124.4]
  wire [31:0] _T_2507; // @[Mux.scala 31:69:@15169.4]
  wire  _T_2484; // @[package.scala 96:25:@15115.4 package.scala 96:25:@15116.4]
  wire [31:0] _T_2508; // @[Mux.scala 31:69:@15170.4]
  wire  _T_2481; // @[package.scala 96:25:@15107.4 package.scala 96:25:@15108.4]
  wire [31:0] _T_2509; // @[Mux.scala 31:69:@15171.4]
  wire  _T_2478; // @[package.scala 96:25:@15099.4 package.scala 96:25:@15100.4]
  wire [31:0] _T_2510; // @[Mux.scala 31:69:@15172.4]
  wire  _T_2475; // @[package.scala 96:25:@15091.4 package.scala 96:25:@15092.4]
  wire [31:0] _T_2511; // @[Mux.scala 31:69:@15173.4]
  wire  _T_2472; // @[package.scala 96:25:@15083.4 package.scala 96:25:@15084.4]
  wire [31:0] _T_2512; // @[Mux.scala 31:69:@15174.4]
  wire  _T_2469; // @[package.scala 96:25:@15075.4 package.scala 96:25:@15076.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12477.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12493.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12509.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12525.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12541.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12557.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12573.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12589.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12605.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12621.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12637.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12653.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@12849.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@12938.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@13027.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13116.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13205.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13294.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13383.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13472.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13561.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13650.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13739.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@13828.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@13918.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@13926.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@13934.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@13942.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@13950.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@13958.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@13966.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@13974.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@13982.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@13990.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@13998.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14006.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14062.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14070.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14078.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14086.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14094.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14102.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14110.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14118.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14126.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14134.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14142.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14150.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14206.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14214.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14222.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14230.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14238.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14246.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14254.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14262.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14270.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14278.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14286.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14294.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14350.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14358.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14366.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14374.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14382.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14390.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14398.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14406.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14414.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14422.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14430.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14438.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14494.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14502.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14510.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14518.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14526.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14534.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14542.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14550.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14558.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14566.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14574.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14582.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14638.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14646.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14654.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14662.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14670.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14678.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14686.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@14694.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@14702.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@14710.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@14718.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@14726.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@14782.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@14790.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@14798.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@14806.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@14814.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@14822.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@14830.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@14838.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@14846.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@14854.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@14862.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@14870.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@14926.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@14934.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@14942.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@14950.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@14958.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@14966.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@14974.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@14982.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@14990.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@14998.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15006.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15014.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@15070.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@15078.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@15086.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@15094.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@15102.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@15110.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@15118.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@15126.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@15134.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@15142.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@15150.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@15158.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  assign _T_316 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12669.4]
  assign _T_318 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@12670.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 82:228:@12671.4]
  assign _T_320 = io_wPort_0_en_0 & _T_319; // @[MemPrimitives.scala 83:102:@12672.4]
  assign _T_322 = {_T_320,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12674.4]
  assign _T_329 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@12682.4]
  assign _T_330 = _T_316 & _T_329; // @[MemPrimitives.scala 82:228:@12683.4]
  assign _T_331 = io_wPort_0_en_0 & _T_330; // @[MemPrimitives.scala 83:102:@12684.4]
  assign _T_333 = {_T_331,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12686.4]
  assign _T_340 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@12694.4]
  assign _T_341 = _T_316 & _T_340; // @[MemPrimitives.scala 82:228:@12695.4]
  assign _T_342 = io_wPort_0_en_0 & _T_341; // @[MemPrimitives.scala 83:102:@12696.4]
  assign _T_344 = {_T_342,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12698.4]
  assign _T_349 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12705.4]
  assign _T_352 = _T_349 & _T_318; // @[MemPrimitives.scala 82:228:@12707.4]
  assign _T_353 = io_wPort_0_en_0 & _T_352; // @[MemPrimitives.scala 83:102:@12708.4]
  assign _T_355 = {_T_353,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12710.4]
  assign _T_363 = _T_349 & _T_329; // @[MemPrimitives.scala 82:228:@12719.4]
  assign _T_364 = io_wPort_0_en_0 & _T_363; // @[MemPrimitives.scala 83:102:@12720.4]
  assign _T_366 = {_T_364,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12722.4]
  assign _T_374 = _T_349 & _T_340; // @[MemPrimitives.scala 82:228:@12731.4]
  assign _T_375 = io_wPort_0_en_0 & _T_374; // @[MemPrimitives.scala 83:102:@12732.4]
  assign _T_377 = {_T_375,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12734.4]
  assign _T_382 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12741.4]
  assign _T_385 = _T_382 & _T_318; // @[MemPrimitives.scala 82:228:@12743.4]
  assign _T_386 = io_wPort_0_en_0 & _T_385; // @[MemPrimitives.scala 83:102:@12744.4]
  assign _T_388 = {_T_386,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12746.4]
  assign _T_396 = _T_382 & _T_329; // @[MemPrimitives.scala 82:228:@12755.4]
  assign _T_397 = io_wPort_0_en_0 & _T_396; // @[MemPrimitives.scala 83:102:@12756.4]
  assign _T_399 = {_T_397,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12758.4]
  assign _T_407 = _T_382 & _T_340; // @[MemPrimitives.scala 82:228:@12767.4]
  assign _T_408 = io_wPort_0_en_0 & _T_407; // @[MemPrimitives.scala 83:102:@12768.4]
  assign _T_410 = {_T_408,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12770.4]
  assign _T_415 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12777.4]
  assign _T_418 = _T_415 & _T_318; // @[MemPrimitives.scala 82:228:@12779.4]
  assign _T_419 = io_wPort_0_en_0 & _T_418; // @[MemPrimitives.scala 83:102:@12780.4]
  assign _T_421 = {_T_419,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12782.4]
  assign _T_429 = _T_415 & _T_329; // @[MemPrimitives.scala 82:228:@12791.4]
  assign _T_430 = io_wPort_0_en_0 & _T_429; // @[MemPrimitives.scala 83:102:@12792.4]
  assign _T_432 = {_T_430,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12794.4]
  assign _T_440 = _T_415 & _T_340; // @[MemPrimitives.scala 82:228:@12803.4]
  assign _T_441 = io_wPort_0_en_0 & _T_440; // @[MemPrimitives.scala 83:102:@12804.4]
  assign _T_443 = {_T_441,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12806.4]
  assign _T_448 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12813.4]
  assign _T_450 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12814.4]
  assign _T_451 = _T_448 & _T_450; // @[MemPrimitives.scala 110:228:@12815.4]
  assign _T_454 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12817.4]
  assign _T_456 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12818.4]
  assign _T_457 = _T_454 & _T_456; // @[MemPrimitives.scala 110:228:@12819.4]
  assign _T_460 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12821.4]
  assign _T_462 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12822.4]
  assign _T_463 = _T_460 & _T_462; // @[MemPrimitives.scala 110:228:@12823.4]
  assign _T_466 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12825.4]
  assign _T_468 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12826.4]
  assign _T_469 = _T_466 & _T_468; // @[MemPrimitives.scala 110:228:@12827.4]
  assign _T_472 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12829.4]
  assign _T_474 = io_rPort_4_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12830.4]
  assign _T_475 = _T_472 & _T_474; // @[MemPrimitives.scala 110:228:@12831.4]
  assign _T_478 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12833.4]
  assign _T_480 = io_rPort_5_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12834.4]
  assign _T_481 = _T_478 & _T_480; // @[MemPrimitives.scala 110:228:@12835.4]
  assign _T_484 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12837.4]
  assign _T_486 = io_rPort_6_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12838.4]
  assign _T_487 = _T_484 & _T_486; // @[MemPrimitives.scala 110:228:@12839.4]
  assign _T_490 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12841.4]
  assign _T_492 = io_rPort_7_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12842.4]
  assign _T_493 = _T_490 & _T_492; // @[MemPrimitives.scala 110:228:@12843.4]
  assign _T_496 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12845.4]
  assign _T_498 = io_rPort_8_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12846.4]
  assign _T_499 = _T_496 & _T_498; // @[MemPrimitives.scala 110:228:@12847.4]
  assign _T_501 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@12861.4]
  assign _T_502 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@12862.4]
  assign _T_503 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@12863.4]
  assign _T_504 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@12864.4]
  assign _T_505 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@12865.4]
  assign _T_506 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@12866.4]
  assign _T_507 = StickySelects_io_outs_6; // @[MemPrimitives.scala 126:35:@12867.4]
  assign _T_508 = StickySelects_io_outs_7; // @[MemPrimitives.scala 126:35:@12868.4]
  assign _T_509 = StickySelects_io_outs_8; // @[MemPrimitives.scala 126:35:@12869.4]
  assign _T_511 = {_T_501,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12871.4]
  assign _T_513 = {_T_502,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12873.4]
  assign _T_515 = {_T_503,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12875.4]
  assign _T_517 = {_T_504,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12877.4]
  assign _T_519 = {_T_505,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12879.4]
  assign _T_521 = {_T_506,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12881.4]
  assign _T_523 = {_T_507,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12883.4]
  assign _T_525 = {_T_508,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12885.4]
  assign _T_527 = {_T_509,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12887.4]
  assign _T_528 = _T_508 ? _T_525 : _T_527; // @[Mux.scala 31:69:@12888.4]
  assign _T_529 = _T_507 ? _T_523 : _T_528; // @[Mux.scala 31:69:@12889.4]
  assign _T_530 = _T_506 ? _T_521 : _T_529; // @[Mux.scala 31:69:@12890.4]
  assign _T_531 = _T_505 ? _T_519 : _T_530; // @[Mux.scala 31:69:@12891.4]
  assign _T_532 = _T_504 ? _T_517 : _T_531; // @[Mux.scala 31:69:@12892.4]
  assign _T_533 = _T_503 ? _T_515 : _T_532; // @[Mux.scala 31:69:@12893.4]
  assign _T_534 = _T_502 ? _T_513 : _T_533; // @[Mux.scala 31:69:@12894.4]
  assign _T_535 = _T_501 ? _T_511 : _T_534; // @[Mux.scala 31:69:@12895.4]
  assign _T_542 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12903.4]
  assign _T_543 = _T_448 & _T_542; // @[MemPrimitives.scala 110:228:@12904.4]
  assign _T_548 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12907.4]
  assign _T_549 = _T_454 & _T_548; // @[MemPrimitives.scala 110:228:@12908.4]
  assign _T_554 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12911.4]
  assign _T_555 = _T_460 & _T_554; // @[MemPrimitives.scala 110:228:@12912.4]
  assign _T_560 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12915.4]
  assign _T_561 = _T_466 & _T_560; // @[MemPrimitives.scala 110:228:@12916.4]
  assign _T_566 = io_rPort_4_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12919.4]
  assign _T_567 = _T_472 & _T_566; // @[MemPrimitives.scala 110:228:@12920.4]
  assign _T_572 = io_rPort_5_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12923.4]
  assign _T_573 = _T_478 & _T_572; // @[MemPrimitives.scala 110:228:@12924.4]
  assign _T_578 = io_rPort_6_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12927.4]
  assign _T_579 = _T_484 & _T_578; // @[MemPrimitives.scala 110:228:@12928.4]
  assign _T_584 = io_rPort_7_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12931.4]
  assign _T_585 = _T_490 & _T_584; // @[MemPrimitives.scala 110:228:@12932.4]
  assign _T_590 = io_rPort_8_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@12935.4]
  assign _T_591 = _T_496 & _T_590; // @[MemPrimitives.scala 110:228:@12936.4]
  assign _T_593 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@12950.4]
  assign _T_594 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@12951.4]
  assign _T_595 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@12952.4]
  assign _T_596 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@12953.4]
  assign _T_597 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@12954.4]
  assign _T_598 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@12955.4]
  assign _T_599 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 126:35:@12956.4]
  assign _T_600 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 126:35:@12957.4]
  assign _T_601 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 126:35:@12958.4]
  assign _T_603 = {_T_593,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12960.4]
  assign _T_605 = {_T_594,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12962.4]
  assign _T_607 = {_T_595,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12964.4]
  assign _T_609 = {_T_596,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12966.4]
  assign _T_611 = {_T_597,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12968.4]
  assign _T_613 = {_T_598,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12970.4]
  assign _T_615 = {_T_599,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12972.4]
  assign _T_617 = {_T_600,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12974.4]
  assign _T_619 = {_T_601,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12976.4]
  assign _T_620 = _T_600 ? _T_617 : _T_619; // @[Mux.scala 31:69:@12977.4]
  assign _T_621 = _T_599 ? _T_615 : _T_620; // @[Mux.scala 31:69:@12978.4]
  assign _T_622 = _T_598 ? _T_613 : _T_621; // @[Mux.scala 31:69:@12979.4]
  assign _T_623 = _T_597 ? _T_611 : _T_622; // @[Mux.scala 31:69:@12980.4]
  assign _T_624 = _T_596 ? _T_609 : _T_623; // @[Mux.scala 31:69:@12981.4]
  assign _T_625 = _T_595 ? _T_607 : _T_624; // @[Mux.scala 31:69:@12982.4]
  assign _T_626 = _T_594 ? _T_605 : _T_625; // @[Mux.scala 31:69:@12983.4]
  assign _T_627 = _T_593 ? _T_603 : _T_626; // @[Mux.scala 31:69:@12984.4]
  assign _T_634 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@12992.4]
  assign _T_635 = _T_448 & _T_634; // @[MemPrimitives.scala 110:228:@12993.4]
  assign _T_640 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@12996.4]
  assign _T_641 = _T_454 & _T_640; // @[MemPrimitives.scala 110:228:@12997.4]
  assign _T_646 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13000.4]
  assign _T_647 = _T_460 & _T_646; // @[MemPrimitives.scala 110:228:@13001.4]
  assign _T_652 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13004.4]
  assign _T_653 = _T_466 & _T_652; // @[MemPrimitives.scala 110:228:@13005.4]
  assign _T_658 = io_rPort_4_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13008.4]
  assign _T_659 = _T_472 & _T_658; // @[MemPrimitives.scala 110:228:@13009.4]
  assign _T_664 = io_rPort_5_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13012.4]
  assign _T_665 = _T_478 & _T_664; // @[MemPrimitives.scala 110:228:@13013.4]
  assign _T_670 = io_rPort_6_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13016.4]
  assign _T_671 = _T_484 & _T_670; // @[MemPrimitives.scala 110:228:@13017.4]
  assign _T_676 = io_rPort_7_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13020.4]
  assign _T_677 = _T_490 & _T_676; // @[MemPrimitives.scala 110:228:@13021.4]
  assign _T_682 = io_rPort_8_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13024.4]
  assign _T_683 = _T_496 & _T_682; // @[MemPrimitives.scala 110:228:@13025.4]
  assign _T_685 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@13039.4]
  assign _T_686 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@13040.4]
  assign _T_687 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@13041.4]
  assign _T_688 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@13042.4]
  assign _T_689 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@13043.4]
  assign _T_690 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@13044.4]
  assign _T_691 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 126:35:@13045.4]
  assign _T_692 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 126:35:@13046.4]
  assign _T_693 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 126:35:@13047.4]
  assign _T_695 = {_T_685,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13049.4]
  assign _T_697 = {_T_686,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13051.4]
  assign _T_699 = {_T_687,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13053.4]
  assign _T_701 = {_T_688,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13055.4]
  assign _T_703 = {_T_689,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13057.4]
  assign _T_705 = {_T_690,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13059.4]
  assign _T_707 = {_T_691,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13061.4]
  assign _T_709 = {_T_692,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13063.4]
  assign _T_711 = {_T_693,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13065.4]
  assign _T_712 = _T_692 ? _T_709 : _T_711; // @[Mux.scala 31:69:@13066.4]
  assign _T_713 = _T_691 ? _T_707 : _T_712; // @[Mux.scala 31:69:@13067.4]
  assign _T_714 = _T_690 ? _T_705 : _T_713; // @[Mux.scala 31:69:@13068.4]
  assign _T_715 = _T_689 ? _T_703 : _T_714; // @[Mux.scala 31:69:@13069.4]
  assign _T_716 = _T_688 ? _T_701 : _T_715; // @[Mux.scala 31:69:@13070.4]
  assign _T_717 = _T_687 ? _T_699 : _T_716; // @[Mux.scala 31:69:@13071.4]
  assign _T_718 = _T_686 ? _T_697 : _T_717; // @[Mux.scala 31:69:@13072.4]
  assign _T_719 = _T_685 ? _T_695 : _T_718; // @[Mux.scala 31:69:@13073.4]
  assign _T_724 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13080.4]
  assign _T_727 = _T_724 & _T_450; // @[MemPrimitives.scala 110:228:@13082.4]
  assign _T_730 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13084.4]
  assign _T_733 = _T_730 & _T_456; // @[MemPrimitives.scala 110:228:@13086.4]
  assign _T_736 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13088.4]
  assign _T_739 = _T_736 & _T_462; // @[MemPrimitives.scala 110:228:@13090.4]
  assign _T_742 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13092.4]
  assign _T_745 = _T_742 & _T_468; // @[MemPrimitives.scala 110:228:@13094.4]
  assign _T_748 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13096.4]
  assign _T_751 = _T_748 & _T_474; // @[MemPrimitives.scala 110:228:@13098.4]
  assign _T_754 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13100.4]
  assign _T_757 = _T_754 & _T_480; // @[MemPrimitives.scala 110:228:@13102.4]
  assign _T_760 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13104.4]
  assign _T_763 = _T_760 & _T_486; // @[MemPrimitives.scala 110:228:@13106.4]
  assign _T_766 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13108.4]
  assign _T_769 = _T_766 & _T_492; // @[MemPrimitives.scala 110:228:@13110.4]
  assign _T_772 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13112.4]
  assign _T_775 = _T_772 & _T_498; // @[MemPrimitives.scala 110:228:@13114.4]
  assign _T_777 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13128.4]
  assign _T_778 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13129.4]
  assign _T_779 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13130.4]
  assign _T_780 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13131.4]
  assign _T_781 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13132.4]
  assign _T_782 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13133.4]
  assign _T_783 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 126:35:@13134.4]
  assign _T_784 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 126:35:@13135.4]
  assign _T_785 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 126:35:@13136.4]
  assign _T_787 = {_T_777,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13138.4]
  assign _T_789 = {_T_778,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13140.4]
  assign _T_791 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13142.4]
  assign _T_793 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13144.4]
  assign _T_795 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13146.4]
  assign _T_797 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13148.4]
  assign _T_799 = {_T_783,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13150.4]
  assign _T_801 = {_T_784,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13152.4]
  assign _T_803 = {_T_785,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13154.4]
  assign _T_804 = _T_784 ? _T_801 : _T_803; // @[Mux.scala 31:69:@13155.4]
  assign _T_805 = _T_783 ? _T_799 : _T_804; // @[Mux.scala 31:69:@13156.4]
  assign _T_806 = _T_782 ? _T_797 : _T_805; // @[Mux.scala 31:69:@13157.4]
  assign _T_807 = _T_781 ? _T_795 : _T_806; // @[Mux.scala 31:69:@13158.4]
  assign _T_808 = _T_780 ? _T_793 : _T_807; // @[Mux.scala 31:69:@13159.4]
  assign _T_809 = _T_779 ? _T_791 : _T_808; // @[Mux.scala 31:69:@13160.4]
  assign _T_810 = _T_778 ? _T_789 : _T_809; // @[Mux.scala 31:69:@13161.4]
  assign _T_811 = _T_777 ? _T_787 : _T_810; // @[Mux.scala 31:69:@13162.4]
  assign _T_819 = _T_724 & _T_542; // @[MemPrimitives.scala 110:228:@13171.4]
  assign _T_825 = _T_730 & _T_548; // @[MemPrimitives.scala 110:228:@13175.4]
  assign _T_831 = _T_736 & _T_554; // @[MemPrimitives.scala 110:228:@13179.4]
  assign _T_837 = _T_742 & _T_560; // @[MemPrimitives.scala 110:228:@13183.4]
  assign _T_843 = _T_748 & _T_566; // @[MemPrimitives.scala 110:228:@13187.4]
  assign _T_849 = _T_754 & _T_572; // @[MemPrimitives.scala 110:228:@13191.4]
  assign _T_855 = _T_760 & _T_578; // @[MemPrimitives.scala 110:228:@13195.4]
  assign _T_861 = _T_766 & _T_584; // @[MemPrimitives.scala 110:228:@13199.4]
  assign _T_867 = _T_772 & _T_590; // @[MemPrimitives.scala 110:228:@13203.4]
  assign _T_869 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13217.4]
  assign _T_870 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13218.4]
  assign _T_871 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13219.4]
  assign _T_872 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13220.4]
  assign _T_873 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13221.4]
  assign _T_874 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13222.4]
  assign _T_875 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 126:35:@13223.4]
  assign _T_876 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 126:35:@13224.4]
  assign _T_877 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 126:35:@13225.4]
  assign _T_879 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13227.4]
  assign _T_881 = {_T_870,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13229.4]
  assign _T_883 = {_T_871,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13231.4]
  assign _T_885 = {_T_872,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13233.4]
  assign _T_887 = {_T_873,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13235.4]
  assign _T_889 = {_T_874,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13237.4]
  assign _T_891 = {_T_875,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13239.4]
  assign _T_893 = {_T_876,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13241.4]
  assign _T_895 = {_T_877,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13243.4]
  assign _T_896 = _T_876 ? _T_893 : _T_895; // @[Mux.scala 31:69:@13244.4]
  assign _T_897 = _T_875 ? _T_891 : _T_896; // @[Mux.scala 31:69:@13245.4]
  assign _T_898 = _T_874 ? _T_889 : _T_897; // @[Mux.scala 31:69:@13246.4]
  assign _T_899 = _T_873 ? _T_887 : _T_898; // @[Mux.scala 31:69:@13247.4]
  assign _T_900 = _T_872 ? _T_885 : _T_899; // @[Mux.scala 31:69:@13248.4]
  assign _T_901 = _T_871 ? _T_883 : _T_900; // @[Mux.scala 31:69:@13249.4]
  assign _T_902 = _T_870 ? _T_881 : _T_901; // @[Mux.scala 31:69:@13250.4]
  assign _T_903 = _T_869 ? _T_879 : _T_902; // @[Mux.scala 31:69:@13251.4]
  assign _T_911 = _T_724 & _T_634; // @[MemPrimitives.scala 110:228:@13260.4]
  assign _T_917 = _T_730 & _T_640; // @[MemPrimitives.scala 110:228:@13264.4]
  assign _T_923 = _T_736 & _T_646; // @[MemPrimitives.scala 110:228:@13268.4]
  assign _T_929 = _T_742 & _T_652; // @[MemPrimitives.scala 110:228:@13272.4]
  assign _T_935 = _T_748 & _T_658; // @[MemPrimitives.scala 110:228:@13276.4]
  assign _T_941 = _T_754 & _T_664; // @[MemPrimitives.scala 110:228:@13280.4]
  assign _T_947 = _T_760 & _T_670; // @[MemPrimitives.scala 110:228:@13284.4]
  assign _T_953 = _T_766 & _T_676; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_959 = _T_772 & _T_682; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_961 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13306.4]
  assign _T_962 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13307.4]
  assign _T_963 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13308.4]
  assign _T_964 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13309.4]
  assign _T_965 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13310.4]
  assign _T_966 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13311.4]
  assign _T_967 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 126:35:@13312.4]
  assign _T_968 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 126:35:@13313.4]
  assign _T_969 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 126:35:@13314.4]
  assign _T_971 = {_T_961,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13316.4]
  assign _T_973 = {_T_962,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13318.4]
  assign _T_975 = {_T_963,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13320.4]
  assign _T_977 = {_T_964,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13322.4]
  assign _T_979 = {_T_965,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13324.4]
  assign _T_981 = {_T_966,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13326.4]
  assign _T_983 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13328.4]
  assign _T_985 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13330.4]
  assign _T_987 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13332.4]
  assign _T_988 = _T_968 ? _T_985 : _T_987; // @[Mux.scala 31:69:@13333.4]
  assign _T_989 = _T_967 ? _T_983 : _T_988; // @[Mux.scala 31:69:@13334.4]
  assign _T_990 = _T_966 ? _T_981 : _T_989; // @[Mux.scala 31:69:@13335.4]
  assign _T_991 = _T_965 ? _T_979 : _T_990; // @[Mux.scala 31:69:@13336.4]
  assign _T_992 = _T_964 ? _T_977 : _T_991; // @[Mux.scala 31:69:@13337.4]
  assign _T_993 = _T_963 ? _T_975 : _T_992; // @[Mux.scala 31:69:@13338.4]
  assign _T_994 = _T_962 ? _T_973 : _T_993; // @[Mux.scala 31:69:@13339.4]
  assign _T_995 = _T_961 ? _T_971 : _T_994; // @[Mux.scala 31:69:@13340.4]
  assign _T_1000 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13347.4]
  assign _T_1003 = _T_1000 & _T_450; // @[MemPrimitives.scala 110:228:@13349.4]
  assign _T_1006 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13351.4]
  assign _T_1009 = _T_1006 & _T_456; // @[MemPrimitives.scala 110:228:@13353.4]
  assign _T_1012 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13355.4]
  assign _T_1015 = _T_1012 & _T_462; // @[MemPrimitives.scala 110:228:@13357.4]
  assign _T_1018 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13359.4]
  assign _T_1021 = _T_1018 & _T_468; // @[MemPrimitives.scala 110:228:@13361.4]
  assign _T_1024 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13363.4]
  assign _T_1027 = _T_1024 & _T_474; // @[MemPrimitives.scala 110:228:@13365.4]
  assign _T_1030 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13367.4]
  assign _T_1033 = _T_1030 & _T_480; // @[MemPrimitives.scala 110:228:@13369.4]
  assign _T_1036 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13371.4]
  assign _T_1039 = _T_1036 & _T_486; // @[MemPrimitives.scala 110:228:@13373.4]
  assign _T_1042 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13375.4]
  assign _T_1045 = _T_1042 & _T_492; // @[MemPrimitives.scala 110:228:@13377.4]
  assign _T_1048 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13379.4]
  assign _T_1051 = _T_1048 & _T_498; // @[MemPrimitives.scala 110:228:@13381.4]
  assign _T_1053 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13395.4]
  assign _T_1054 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13396.4]
  assign _T_1055 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13397.4]
  assign _T_1056 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13398.4]
  assign _T_1057 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13399.4]
  assign _T_1058 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13400.4]
  assign _T_1059 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 126:35:@13401.4]
  assign _T_1060 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 126:35:@13402.4]
  assign _T_1061 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 126:35:@13403.4]
  assign _T_1063 = {_T_1053,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13405.4]
  assign _T_1065 = {_T_1054,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13407.4]
  assign _T_1067 = {_T_1055,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13409.4]
  assign _T_1069 = {_T_1056,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13411.4]
  assign _T_1071 = {_T_1057,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13413.4]
  assign _T_1073 = {_T_1058,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13415.4]
  assign _T_1075 = {_T_1059,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13417.4]
  assign _T_1077 = {_T_1060,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13419.4]
  assign _T_1079 = {_T_1061,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13421.4]
  assign _T_1080 = _T_1060 ? _T_1077 : _T_1079; // @[Mux.scala 31:69:@13422.4]
  assign _T_1081 = _T_1059 ? _T_1075 : _T_1080; // @[Mux.scala 31:69:@13423.4]
  assign _T_1082 = _T_1058 ? _T_1073 : _T_1081; // @[Mux.scala 31:69:@13424.4]
  assign _T_1083 = _T_1057 ? _T_1071 : _T_1082; // @[Mux.scala 31:69:@13425.4]
  assign _T_1084 = _T_1056 ? _T_1069 : _T_1083; // @[Mux.scala 31:69:@13426.4]
  assign _T_1085 = _T_1055 ? _T_1067 : _T_1084; // @[Mux.scala 31:69:@13427.4]
  assign _T_1086 = _T_1054 ? _T_1065 : _T_1085; // @[Mux.scala 31:69:@13428.4]
  assign _T_1087 = _T_1053 ? _T_1063 : _T_1086; // @[Mux.scala 31:69:@13429.4]
  assign _T_1095 = _T_1000 & _T_542; // @[MemPrimitives.scala 110:228:@13438.4]
  assign _T_1101 = _T_1006 & _T_548; // @[MemPrimitives.scala 110:228:@13442.4]
  assign _T_1107 = _T_1012 & _T_554; // @[MemPrimitives.scala 110:228:@13446.4]
  assign _T_1113 = _T_1018 & _T_560; // @[MemPrimitives.scala 110:228:@13450.4]
  assign _T_1119 = _T_1024 & _T_566; // @[MemPrimitives.scala 110:228:@13454.4]
  assign _T_1125 = _T_1030 & _T_572; // @[MemPrimitives.scala 110:228:@13458.4]
  assign _T_1131 = _T_1036 & _T_578; // @[MemPrimitives.scala 110:228:@13462.4]
  assign _T_1137 = _T_1042 & _T_584; // @[MemPrimitives.scala 110:228:@13466.4]
  assign _T_1143 = _T_1048 & _T_590; // @[MemPrimitives.scala 110:228:@13470.4]
  assign _T_1145 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13484.4]
  assign _T_1146 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13485.4]
  assign _T_1147 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13486.4]
  assign _T_1148 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13487.4]
  assign _T_1149 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13488.4]
  assign _T_1150 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13489.4]
  assign _T_1151 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 126:35:@13490.4]
  assign _T_1152 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 126:35:@13491.4]
  assign _T_1153 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 126:35:@13492.4]
  assign _T_1155 = {_T_1145,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13494.4]
  assign _T_1157 = {_T_1146,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13496.4]
  assign _T_1159 = {_T_1147,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13498.4]
  assign _T_1161 = {_T_1148,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13500.4]
  assign _T_1163 = {_T_1149,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13502.4]
  assign _T_1165 = {_T_1150,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13504.4]
  assign _T_1167 = {_T_1151,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13506.4]
  assign _T_1169 = {_T_1152,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13508.4]
  assign _T_1171 = {_T_1153,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13510.4]
  assign _T_1172 = _T_1152 ? _T_1169 : _T_1171; // @[Mux.scala 31:69:@13511.4]
  assign _T_1173 = _T_1151 ? _T_1167 : _T_1172; // @[Mux.scala 31:69:@13512.4]
  assign _T_1174 = _T_1150 ? _T_1165 : _T_1173; // @[Mux.scala 31:69:@13513.4]
  assign _T_1175 = _T_1149 ? _T_1163 : _T_1174; // @[Mux.scala 31:69:@13514.4]
  assign _T_1176 = _T_1148 ? _T_1161 : _T_1175; // @[Mux.scala 31:69:@13515.4]
  assign _T_1177 = _T_1147 ? _T_1159 : _T_1176; // @[Mux.scala 31:69:@13516.4]
  assign _T_1178 = _T_1146 ? _T_1157 : _T_1177; // @[Mux.scala 31:69:@13517.4]
  assign _T_1179 = _T_1145 ? _T_1155 : _T_1178; // @[Mux.scala 31:69:@13518.4]
  assign _T_1187 = _T_1000 & _T_634; // @[MemPrimitives.scala 110:228:@13527.4]
  assign _T_1193 = _T_1006 & _T_640; // @[MemPrimitives.scala 110:228:@13531.4]
  assign _T_1199 = _T_1012 & _T_646; // @[MemPrimitives.scala 110:228:@13535.4]
  assign _T_1205 = _T_1018 & _T_652; // @[MemPrimitives.scala 110:228:@13539.4]
  assign _T_1211 = _T_1024 & _T_658; // @[MemPrimitives.scala 110:228:@13543.4]
  assign _T_1217 = _T_1030 & _T_664; // @[MemPrimitives.scala 110:228:@13547.4]
  assign _T_1223 = _T_1036 & _T_670; // @[MemPrimitives.scala 110:228:@13551.4]
  assign _T_1229 = _T_1042 & _T_676; // @[MemPrimitives.scala 110:228:@13555.4]
  assign _T_1235 = _T_1048 & _T_682; // @[MemPrimitives.scala 110:228:@13559.4]
  assign _T_1237 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13573.4]
  assign _T_1238 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13574.4]
  assign _T_1239 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13575.4]
  assign _T_1240 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13576.4]
  assign _T_1241 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13577.4]
  assign _T_1242 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13578.4]
  assign _T_1243 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 126:35:@13579.4]
  assign _T_1244 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 126:35:@13580.4]
  assign _T_1245 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 126:35:@13581.4]
  assign _T_1247 = {_T_1237,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13583.4]
  assign _T_1249 = {_T_1238,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13585.4]
  assign _T_1251 = {_T_1239,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13587.4]
  assign _T_1253 = {_T_1240,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13589.4]
  assign _T_1255 = {_T_1241,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13591.4]
  assign _T_1257 = {_T_1242,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13593.4]
  assign _T_1259 = {_T_1243,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13595.4]
  assign _T_1261 = {_T_1244,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13597.4]
  assign _T_1263 = {_T_1245,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13599.4]
  assign _T_1264 = _T_1244 ? _T_1261 : _T_1263; // @[Mux.scala 31:69:@13600.4]
  assign _T_1265 = _T_1243 ? _T_1259 : _T_1264; // @[Mux.scala 31:69:@13601.4]
  assign _T_1266 = _T_1242 ? _T_1257 : _T_1265; // @[Mux.scala 31:69:@13602.4]
  assign _T_1267 = _T_1241 ? _T_1255 : _T_1266; // @[Mux.scala 31:69:@13603.4]
  assign _T_1268 = _T_1240 ? _T_1253 : _T_1267; // @[Mux.scala 31:69:@13604.4]
  assign _T_1269 = _T_1239 ? _T_1251 : _T_1268; // @[Mux.scala 31:69:@13605.4]
  assign _T_1270 = _T_1238 ? _T_1249 : _T_1269; // @[Mux.scala 31:69:@13606.4]
  assign _T_1271 = _T_1237 ? _T_1247 : _T_1270; // @[Mux.scala 31:69:@13607.4]
  assign _T_1276 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13614.4]
  assign _T_1279 = _T_1276 & _T_450; // @[MemPrimitives.scala 110:228:@13616.4]
  assign _T_1282 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13618.4]
  assign _T_1285 = _T_1282 & _T_456; // @[MemPrimitives.scala 110:228:@13620.4]
  assign _T_1288 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13622.4]
  assign _T_1291 = _T_1288 & _T_462; // @[MemPrimitives.scala 110:228:@13624.4]
  assign _T_1294 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13626.4]
  assign _T_1297 = _T_1294 & _T_468; // @[MemPrimitives.scala 110:228:@13628.4]
  assign _T_1300 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13630.4]
  assign _T_1303 = _T_1300 & _T_474; // @[MemPrimitives.scala 110:228:@13632.4]
  assign _T_1306 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13634.4]
  assign _T_1309 = _T_1306 & _T_480; // @[MemPrimitives.scala 110:228:@13636.4]
  assign _T_1312 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13638.4]
  assign _T_1315 = _T_1312 & _T_486; // @[MemPrimitives.scala 110:228:@13640.4]
  assign _T_1318 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13642.4]
  assign _T_1321 = _T_1318 & _T_492; // @[MemPrimitives.scala 110:228:@13644.4]
  assign _T_1324 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13646.4]
  assign _T_1327 = _T_1324 & _T_498; // @[MemPrimitives.scala 110:228:@13648.4]
  assign _T_1329 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13662.4]
  assign _T_1330 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13663.4]
  assign _T_1331 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13664.4]
  assign _T_1332 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13665.4]
  assign _T_1333 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13666.4]
  assign _T_1334 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13667.4]
  assign _T_1335 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 126:35:@13668.4]
  assign _T_1336 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 126:35:@13669.4]
  assign _T_1337 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 126:35:@13670.4]
  assign _T_1339 = {_T_1329,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13672.4]
  assign _T_1341 = {_T_1330,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13674.4]
  assign _T_1343 = {_T_1331,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13676.4]
  assign _T_1345 = {_T_1332,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13678.4]
  assign _T_1347 = {_T_1333,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13680.4]
  assign _T_1349 = {_T_1334,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13682.4]
  assign _T_1351 = {_T_1335,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13684.4]
  assign _T_1353 = {_T_1336,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13686.4]
  assign _T_1355 = {_T_1337,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13688.4]
  assign _T_1356 = _T_1336 ? _T_1353 : _T_1355; // @[Mux.scala 31:69:@13689.4]
  assign _T_1357 = _T_1335 ? _T_1351 : _T_1356; // @[Mux.scala 31:69:@13690.4]
  assign _T_1358 = _T_1334 ? _T_1349 : _T_1357; // @[Mux.scala 31:69:@13691.4]
  assign _T_1359 = _T_1333 ? _T_1347 : _T_1358; // @[Mux.scala 31:69:@13692.4]
  assign _T_1360 = _T_1332 ? _T_1345 : _T_1359; // @[Mux.scala 31:69:@13693.4]
  assign _T_1361 = _T_1331 ? _T_1343 : _T_1360; // @[Mux.scala 31:69:@13694.4]
  assign _T_1362 = _T_1330 ? _T_1341 : _T_1361; // @[Mux.scala 31:69:@13695.4]
  assign _T_1363 = _T_1329 ? _T_1339 : _T_1362; // @[Mux.scala 31:69:@13696.4]
  assign _T_1371 = _T_1276 & _T_542; // @[MemPrimitives.scala 110:228:@13705.4]
  assign _T_1377 = _T_1282 & _T_548; // @[MemPrimitives.scala 110:228:@13709.4]
  assign _T_1383 = _T_1288 & _T_554; // @[MemPrimitives.scala 110:228:@13713.4]
  assign _T_1389 = _T_1294 & _T_560; // @[MemPrimitives.scala 110:228:@13717.4]
  assign _T_1395 = _T_1300 & _T_566; // @[MemPrimitives.scala 110:228:@13721.4]
  assign _T_1401 = _T_1306 & _T_572; // @[MemPrimitives.scala 110:228:@13725.4]
  assign _T_1407 = _T_1312 & _T_578; // @[MemPrimitives.scala 110:228:@13729.4]
  assign _T_1413 = _T_1318 & _T_584; // @[MemPrimitives.scala 110:228:@13733.4]
  assign _T_1419 = _T_1324 & _T_590; // @[MemPrimitives.scala 110:228:@13737.4]
  assign _T_1421 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13751.4]
  assign _T_1422 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13752.4]
  assign _T_1423 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13753.4]
  assign _T_1424 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13754.4]
  assign _T_1425 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13755.4]
  assign _T_1426 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13756.4]
  assign _T_1427 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 126:35:@13757.4]
  assign _T_1428 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 126:35:@13758.4]
  assign _T_1429 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 126:35:@13759.4]
  assign _T_1431 = {_T_1421,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13761.4]
  assign _T_1433 = {_T_1422,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13763.4]
  assign _T_1435 = {_T_1423,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13765.4]
  assign _T_1437 = {_T_1424,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13767.4]
  assign _T_1439 = {_T_1425,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13769.4]
  assign _T_1441 = {_T_1426,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13771.4]
  assign _T_1443 = {_T_1427,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13773.4]
  assign _T_1445 = {_T_1428,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13775.4]
  assign _T_1447 = {_T_1429,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13777.4]
  assign _T_1448 = _T_1428 ? _T_1445 : _T_1447; // @[Mux.scala 31:69:@13778.4]
  assign _T_1449 = _T_1427 ? _T_1443 : _T_1448; // @[Mux.scala 31:69:@13779.4]
  assign _T_1450 = _T_1426 ? _T_1441 : _T_1449; // @[Mux.scala 31:69:@13780.4]
  assign _T_1451 = _T_1425 ? _T_1439 : _T_1450; // @[Mux.scala 31:69:@13781.4]
  assign _T_1452 = _T_1424 ? _T_1437 : _T_1451; // @[Mux.scala 31:69:@13782.4]
  assign _T_1453 = _T_1423 ? _T_1435 : _T_1452; // @[Mux.scala 31:69:@13783.4]
  assign _T_1454 = _T_1422 ? _T_1433 : _T_1453; // @[Mux.scala 31:69:@13784.4]
  assign _T_1455 = _T_1421 ? _T_1431 : _T_1454; // @[Mux.scala 31:69:@13785.4]
  assign _T_1463 = _T_1276 & _T_634; // @[MemPrimitives.scala 110:228:@13794.4]
  assign _T_1469 = _T_1282 & _T_640; // @[MemPrimitives.scala 110:228:@13798.4]
  assign _T_1475 = _T_1288 & _T_646; // @[MemPrimitives.scala 110:228:@13802.4]
  assign _T_1481 = _T_1294 & _T_652; // @[MemPrimitives.scala 110:228:@13806.4]
  assign _T_1487 = _T_1300 & _T_658; // @[MemPrimitives.scala 110:228:@13810.4]
  assign _T_1493 = _T_1306 & _T_664; // @[MemPrimitives.scala 110:228:@13814.4]
  assign _T_1499 = _T_1312 & _T_670; // @[MemPrimitives.scala 110:228:@13818.4]
  assign _T_1505 = _T_1318 & _T_676; // @[MemPrimitives.scala 110:228:@13822.4]
  assign _T_1511 = _T_1324 & _T_682; // @[MemPrimitives.scala 110:228:@13826.4]
  assign _T_1513 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@13840.4]
  assign _T_1514 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@13841.4]
  assign _T_1515 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@13842.4]
  assign _T_1516 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@13843.4]
  assign _T_1517 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@13844.4]
  assign _T_1518 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@13845.4]
  assign _T_1519 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 126:35:@13846.4]
  assign _T_1520 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 126:35:@13847.4]
  assign _T_1521 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 126:35:@13848.4]
  assign _T_1523 = {_T_1513,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13850.4]
  assign _T_1525 = {_T_1514,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13852.4]
  assign _T_1527 = {_T_1515,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13854.4]
  assign _T_1529 = {_T_1516,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13856.4]
  assign _T_1531 = {_T_1517,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13858.4]
  assign _T_1533 = {_T_1518,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13860.4]
  assign _T_1535 = {_T_1519,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13862.4]
  assign _T_1537 = {_T_1520,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13864.4]
  assign _T_1539 = {_T_1521,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13866.4]
  assign _T_1540 = _T_1520 ? _T_1537 : _T_1539; // @[Mux.scala 31:69:@13867.4]
  assign _T_1541 = _T_1519 ? _T_1535 : _T_1540; // @[Mux.scala 31:69:@13868.4]
  assign _T_1542 = _T_1518 ? _T_1533 : _T_1541; // @[Mux.scala 31:69:@13869.4]
  assign _T_1543 = _T_1517 ? _T_1531 : _T_1542; // @[Mux.scala 31:69:@13870.4]
  assign _T_1544 = _T_1516 ? _T_1529 : _T_1543; // @[Mux.scala 31:69:@13871.4]
  assign _T_1545 = _T_1515 ? _T_1527 : _T_1544; // @[Mux.scala 31:69:@13872.4]
  assign _T_1546 = _T_1514 ? _T_1525 : _T_1545; // @[Mux.scala 31:69:@13873.4]
  assign _T_1547 = _T_1513 ? _T_1523 : _T_1546; // @[Mux.scala 31:69:@13874.4]
  assign _T_1643 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14003.4 package.scala 96:25:@14004.4]
  assign _T_1647 = _T_1643 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14013.4]
  assign _T_1640 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@13995.4 package.scala 96:25:@13996.4]
  assign _T_1648 = _T_1640 ? Mem1D_9_io_output : _T_1647; // @[Mux.scala 31:69:@14014.4]
  assign _T_1637 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@13987.4 package.scala 96:25:@13988.4]
  assign _T_1649 = _T_1637 ? Mem1D_8_io_output : _T_1648; // @[Mux.scala 31:69:@14015.4]
  assign _T_1634 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@13979.4 package.scala 96:25:@13980.4]
  assign _T_1650 = _T_1634 ? Mem1D_7_io_output : _T_1649; // @[Mux.scala 31:69:@14016.4]
  assign _T_1631 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@13971.4 package.scala 96:25:@13972.4]
  assign _T_1651 = _T_1631 ? Mem1D_6_io_output : _T_1650; // @[Mux.scala 31:69:@14017.4]
  assign _T_1628 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@13963.4 package.scala 96:25:@13964.4]
  assign _T_1652 = _T_1628 ? Mem1D_5_io_output : _T_1651; // @[Mux.scala 31:69:@14018.4]
  assign _T_1625 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@13955.4 package.scala 96:25:@13956.4]
  assign _T_1653 = _T_1625 ? Mem1D_4_io_output : _T_1652; // @[Mux.scala 31:69:@14019.4]
  assign _T_1622 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@13947.4 package.scala 96:25:@13948.4]
  assign _T_1654 = _T_1622 ? Mem1D_3_io_output : _T_1653; // @[Mux.scala 31:69:@14020.4]
  assign _T_1619 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@13939.4 package.scala 96:25:@13940.4]
  assign _T_1655 = _T_1619 ? Mem1D_2_io_output : _T_1654; // @[Mux.scala 31:69:@14021.4]
  assign _T_1616 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@13931.4 package.scala 96:25:@13932.4]
  assign _T_1656 = _T_1616 ? Mem1D_1_io_output : _T_1655; // @[Mux.scala 31:69:@14022.4]
  assign _T_1613 = RetimeWrapper_io_out; // @[package.scala 96:25:@13923.4 package.scala 96:25:@13924.4]
  assign _T_1750 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14147.4 package.scala 96:25:@14148.4]
  assign _T_1754 = _T_1750 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14157.4]
  assign _T_1747 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14139.4 package.scala 96:25:@14140.4]
  assign _T_1755 = _T_1747 ? Mem1D_9_io_output : _T_1754; // @[Mux.scala 31:69:@14158.4]
  assign _T_1744 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14131.4 package.scala 96:25:@14132.4]
  assign _T_1756 = _T_1744 ? Mem1D_8_io_output : _T_1755; // @[Mux.scala 31:69:@14159.4]
  assign _T_1741 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14123.4 package.scala 96:25:@14124.4]
  assign _T_1757 = _T_1741 ? Mem1D_7_io_output : _T_1756; // @[Mux.scala 31:69:@14160.4]
  assign _T_1738 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14115.4 package.scala 96:25:@14116.4]
  assign _T_1758 = _T_1738 ? Mem1D_6_io_output : _T_1757; // @[Mux.scala 31:69:@14161.4]
  assign _T_1735 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14107.4 package.scala 96:25:@14108.4]
  assign _T_1759 = _T_1735 ? Mem1D_5_io_output : _T_1758; // @[Mux.scala 31:69:@14162.4]
  assign _T_1732 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14099.4 package.scala 96:25:@14100.4]
  assign _T_1760 = _T_1732 ? Mem1D_4_io_output : _T_1759; // @[Mux.scala 31:69:@14163.4]
  assign _T_1729 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@14091.4 package.scala 96:25:@14092.4]
  assign _T_1761 = _T_1729 ? Mem1D_3_io_output : _T_1760; // @[Mux.scala 31:69:@14164.4]
  assign _T_1726 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14083.4 package.scala 96:25:@14084.4]
  assign _T_1762 = _T_1726 ? Mem1D_2_io_output : _T_1761; // @[Mux.scala 31:69:@14165.4]
  assign _T_1723 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14075.4 package.scala 96:25:@14076.4]
  assign _T_1763 = _T_1723 ? Mem1D_1_io_output : _T_1762; // @[Mux.scala 31:69:@14166.4]
  assign _T_1720 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14067.4 package.scala 96:25:@14068.4]
  assign _T_1857 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14291.4 package.scala 96:25:@14292.4]
  assign _T_1861 = _T_1857 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14301.4]
  assign _T_1854 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14283.4 package.scala 96:25:@14284.4]
  assign _T_1862 = _T_1854 ? Mem1D_9_io_output : _T_1861; // @[Mux.scala 31:69:@14302.4]
  assign _T_1851 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14275.4 package.scala 96:25:@14276.4]
  assign _T_1863 = _T_1851 ? Mem1D_8_io_output : _T_1862; // @[Mux.scala 31:69:@14303.4]
  assign _T_1848 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@14267.4 package.scala 96:25:@14268.4]
  assign _T_1864 = _T_1848 ? Mem1D_7_io_output : _T_1863; // @[Mux.scala 31:69:@14304.4]
  assign _T_1845 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14259.4 package.scala 96:25:@14260.4]
  assign _T_1865 = _T_1845 ? Mem1D_6_io_output : _T_1864; // @[Mux.scala 31:69:@14305.4]
  assign _T_1842 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14251.4 package.scala 96:25:@14252.4]
  assign _T_1866 = _T_1842 ? Mem1D_5_io_output : _T_1865; // @[Mux.scala 31:69:@14306.4]
  assign _T_1839 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14243.4 package.scala 96:25:@14244.4]
  assign _T_1867 = _T_1839 ? Mem1D_4_io_output : _T_1866; // @[Mux.scala 31:69:@14307.4]
  assign _T_1836 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14235.4 package.scala 96:25:@14236.4]
  assign _T_1868 = _T_1836 ? Mem1D_3_io_output : _T_1867; // @[Mux.scala 31:69:@14308.4]
  assign _T_1833 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14227.4 package.scala 96:25:@14228.4]
  assign _T_1869 = _T_1833 ? Mem1D_2_io_output : _T_1868; // @[Mux.scala 31:69:@14309.4]
  assign _T_1830 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14219.4 package.scala 96:25:@14220.4]
  assign _T_1870 = _T_1830 ? Mem1D_1_io_output : _T_1869; // @[Mux.scala 31:69:@14310.4]
  assign _T_1827 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14211.4 package.scala 96:25:@14212.4]
  assign _T_1964 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14435.4 package.scala 96:25:@14436.4]
  assign _T_1968 = _T_1964 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14445.4]
  assign _T_1961 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14427.4 package.scala 96:25:@14428.4]
  assign _T_1969 = _T_1961 ? Mem1D_9_io_output : _T_1968; // @[Mux.scala 31:69:@14446.4]
  assign _T_1958 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14419.4 package.scala 96:25:@14420.4]
  assign _T_1970 = _T_1958 ? Mem1D_8_io_output : _T_1969; // @[Mux.scala 31:69:@14447.4]
  assign _T_1955 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14411.4 package.scala 96:25:@14412.4]
  assign _T_1971 = _T_1955 ? Mem1D_7_io_output : _T_1970; // @[Mux.scala 31:69:@14448.4]
  assign _T_1952 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14403.4 package.scala 96:25:@14404.4]
  assign _T_1972 = _T_1952 ? Mem1D_6_io_output : _T_1971; // @[Mux.scala 31:69:@14449.4]
  assign _T_1949 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14395.4 package.scala 96:25:@14396.4]
  assign _T_1973 = _T_1949 ? Mem1D_5_io_output : _T_1972; // @[Mux.scala 31:69:@14450.4]
  assign _T_1946 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14387.4 package.scala 96:25:@14388.4]
  assign _T_1974 = _T_1946 ? Mem1D_4_io_output : _T_1973; // @[Mux.scala 31:69:@14451.4]
  assign _T_1943 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@14379.4 package.scala 96:25:@14380.4]
  assign _T_1975 = _T_1943 ? Mem1D_3_io_output : _T_1974; // @[Mux.scala 31:69:@14452.4]
  assign _T_1940 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14371.4 package.scala 96:25:@14372.4]
  assign _T_1976 = _T_1940 ? Mem1D_2_io_output : _T_1975; // @[Mux.scala 31:69:@14453.4]
  assign _T_1937 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14363.4 package.scala 96:25:@14364.4]
  assign _T_1977 = _T_1937 ? Mem1D_1_io_output : _T_1976; // @[Mux.scala 31:69:@14454.4]
  assign _T_1934 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14355.4 package.scala 96:25:@14356.4]
  assign _T_2071 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14579.4 package.scala 96:25:@14580.4]
  assign _T_2075 = _T_2071 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14589.4]
  assign _T_2068 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14571.4 package.scala 96:25:@14572.4]
  assign _T_2076 = _T_2068 ? Mem1D_9_io_output : _T_2075; // @[Mux.scala 31:69:@14590.4]
  assign _T_2065 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14563.4 package.scala 96:25:@14564.4]
  assign _T_2077 = _T_2065 ? Mem1D_8_io_output : _T_2076; // @[Mux.scala 31:69:@14591.4]
  assign _T_2062 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@14555.4 package.scala 96:25:@14556.4]
  assign _T_2078 = _T_2062 ? Mem1D_7_io_output : _T_2077; // @[Mux.scala 31:69:@14592.4]
  assign _T_2059 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14547.4 package.scala 96:25:@14548.4]
  assign _T_2079 = _T_2059 ? Mem1D_6_io_output : _T_2078; // @[Mux.scala 31:69:@14593.4]
  assign _T_2056 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14539.4 package.scala 96:25:@14540.4]
  assign _T_2080 = _T_2056 ? Mem1D_5_io_output : _T_2079; // @[Mux.scala 31:69:@14594.4]
  assign _T_2053 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14531.4 package.scala 96:25:@14532.4]
  assign _T_2081 = _T_2053 ? Mem1D_4_io_output : _T_2080; // @[Mux.scala 31:69:@14595.4]
  assign _T_2050 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14523.4 package.scala 96:25:@14524.4]
  assign _T_2082 = _T_2050 ? Mem1D_3_io_output : _T_2081; // @[Mux.scala 31:69:@14596.4]
  assign _T_2047 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14515.4 package.scala 96:25:@14516.4]
  assign _T_2083 = _T_2047 ? Mem1D_2_io_output : _T_2082; // @[Mux.scala 31:69:@14597.4]
  assign _T_2044 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14507.4 package.scala 96:25:@14508.4]
  assign _T_2084 = _T_2044 ? Mem1D_1_io_output : _T_2083; // @[Mux.scala 31:69:@14598.4]
  assign _T_2041 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14499.4 package.scala 96:25:@14500.4]
  assign _T_2178 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14723.4 package.scala 96:25:@14724.4]
  assign _T_2182 = _T_2178 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14733.4]
  assign _T_2175 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14715.4 package.scala 96:25:@14716.4]
  assign _T_2183 = _T_2175 ? Mem1D_9_io_output : _T_2182; // @[Mux.scala 31:69:@14734.4]
  assign _T_2172 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14707.4 package.scala 96:25:@14708.4]
  assign _T_2184 = _T_2172 ? Mem1D_8_io_output : _T_2183; // @[Mux.scala 31:69:@14735.4]
  assign _T_2169 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14699.4 package.scala 96:25:@14700.4]
  assign _T_2185 = _T_2169 ? Mem1D_7_io_output : _T_2184; // @[Mux.scala 31:69:@14736.4]
  assign _T_2166 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14691.4 package.scala 96:25:@14692.4]
  assign _T_2186 = _T_2166 ? Mem1D_6_io_output : _T_2185; // @[Mux.scala 31:69:@14737.4]
  assign _T_2163 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14683.4 package.scala 96:25:@14684.4]
  assign _T_2187 = _T_2163 ? Mem1D_5_io_output : _T_2186; // @[Mux.scala 31:69:@14738.4]
  assign _T_2160 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14675.4 package.scala 96:25:@14676.4]
  assign _T_2188 = _T_2160 ? Mem1D_4_io_output : _T_2187; // @[Mux.scala 31:69:@14739.4]
  assign _T_2157 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@14667.4 package.scala 96:25:@14668.4]
  assign _T_2189 = _T_2157 ? Mem1D_3_io_output : _T_2188; // @[Mux.scala 31:69:@14740.4]
  assign _T_2154 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14659.4 package.scala 96:25:@14660.4]
  assign _T_2190 = _T_2154 ? Mem1D_2_io_output : _T_2189; // @[Mux.scala 31:69:@14741.4]
  assign _T_2151 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14651.4 package.scala 96:25:@14652.4]
  assign _T_2191 = _T_2151 ? Mem1D_1_io_output : _T_2190; // @[Mux.scala 31:69:@14742.4]
  assign _T_2148 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14643.4 package.scala 96:25:@14644.4]
  assign _T_2285 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@14867.4 package.scala 96:25:@14868.4]
  assign _T_2289 = _T_2285 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14877.4]
  assign _T_2282 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@14859.4 package.scala 96:25:@14860.4]
  assign _T_2290 = _T_2282 ? Mem1D_9_io_output : _T_2289; // @[Mux.scala 31:69:@14878.4]
  assign _T_2279 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@14851.4 package.scala 96:25:@14852.4]
  assign _T_2291 = _T_2279 ? Mem1D_8_io_output : _T_2290; // @[Mux.scala 31:69:@14879.4]
  assign _T_2276 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@14843.4 package.scala 96:25:@14844.4]
  assign _T_2292 = _T_2276 ? Mem1D_7_io_output : _T_2291; // @[Mux.scala 31:69:@14880.4]
  assign _T_2273 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@14835.4 package.scala 96:25:@14836.4]
  assign _T_2293 = _T_2273 ? Mem1D_6_io_output : _T_2292; // @[Mux.scala 31:69:@14881.4]
  assign _T_2270 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@14827.4 package.scala 96:25:@14828.4]
  assign _T_2294 = _T_2270 ? Mem1D_5_io_output : _T_2293; // @[Mux.scala 31:69:@14882.4]
  assign _T_2267 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@14819.4 package.scala 96:25:@14820.4]
  assign _T_2295 = _T_2267 ? Mem1D_4_io_output : _T_2294; // @[Mux.scala 31:69:@14883.4]
  assign _T_2264 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@14811.4 package.scala 96:25:@14812.4]
  assign _T_2296 = _T_2264 ? Mem1D_3_io_output : _T_2295; // @[Mux.scala 31:69:@14884.4]
  assign _T_2261 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14803.4 package.scala 96:25:@14804.4]
  assign _T_2297 = _T_2261 ? Mem1D_2_io_output : _T_2296; // @[Mux.scala 31:69:@14885.4]
  assign _T_2258 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14795.4 package.scala 96:25:@14796.4]
  assign _T_2298 = _T_2258 ? Mem1D_1_io_output : _T_2297; // @[Mux.scala 31:69:@14886.4]
  assign _T_2255 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14787.4 package.scala 96:25:@14788.4]
  assign _T_2392 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15011.4 package.scala 96:25:@15012.4]
  assign _T_2396 = _T_2392 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15021.4]
  assign _T_2389 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15003.4 package.scala 96:25:@15004.4]
  assign _T_2397 = _T_2389 ? Mem1D_9_io_output : _T_2396; // @[Mux.scala 31:69:@15022.4]
  assign _T_2386 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@14995.4 package.scala 96:25:@14996.4]
  assign _T_2398 = _T_2386 ? Mem1D_8_io_output : _T_2397; // @[Mux.scala 31:69:@15023.4]
  assign _T_2383 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@14987.4 package.scala 96:25:@14988.4]
  assign _T_2399 = _T_2383 ? Mem1D_7_io_output : _T_2398; // @[Mux.scala 31:69:@15024.4]
  assign _T_2380 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@14979.4 package.scala 96:25:@14980.4]
  assign _T_2400 = _T_2380 ? Mem1D_6_io_output : _T_2399; // @[Mux.scala 31:69:@15025.4]
  assign _T_2377 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@14971.4 package.scala 96:25:@14972.4]
  assign _T_2401 = _T_2377 ? Mem1D_5_io_output : _T_2400; // @[Mux.scala 31:69:@15026.4]
  assign _T_2374 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@14963.4 package.scala 96:25:@14964.4]
  assign _T_2402 = _T_2374 ? Mem1D_4_io_output : _T_2401; // @[Mux.scala 31:69:@15027.4]
  assign _T_2371 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@14955.4 package.scala 96:25:@14956.4]
  assign _T_2403 = _T_2371 ? Mem1D_3_io_output : _T_2402; // @[Mux.scala 31:69:@15028.4]
  assign _T_2368 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@14947.4 package.scala 96:25:@14948.4]
  assign _T_2404 = _T_2368 ? Mem1D_2_io_output : _T_2403; // @[Mux.scala 31:69:@15029.4]
  assign _T_2365 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@14939.4 package.scala 96:25:@14940.4]
  assign _T_2405 = _T_2365 ? Mem1D_1_io_output : _T_2404; // @[Mux.scala 31:69:@15030.4]
  assign _T_2362 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@14931.4 package.scala 96:25:@14932.4]
  assign _T_2499 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@15155.4 package.scala 96:25:@15156.4]
  assign _T_2503 = _T_2499 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15165.4]
  assign _T_2496 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@15147.4 package.scala 96:25:@15148.4]
  assign _T_2504 = _T_2496 ? Mem1D_9_io_output : _T_2503; // @[Mux.scala 31:69:@15166.4]
  assign _T_2493 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@15139.4 package.scala 96:25:@15140.4]
  assign _T_2505 = _T_2493 ? Mem1D_8_io_output : _T_2504; // @[Mux.scala 31:69:@15167.4]
  assign _T_2490 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@15131.4 package.scala 96:25:@15132.4]
  assign _T_2506 = _T_2490 ? Mem1D_7_io_output : _T_2505; // @[Mux.scala 31:69:@15168.4]
  assign _T_2487 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@15123.4 package.scala 96:25:@15124.4]
  assign _T_2507 = _T_2487 ? Mem1D_6_io_output : _T_2506; // @[Mux.scala 31:69:@15169.4]
  assign _T_2484 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@15115.4 package.scala 96:25:@15116.4]
  assign _T_2508 = _T_2484 ? Mem1D_5_io_output : _T_2507; // @[Mux.scala 31:69:@15170.4]
  assign _T_2481 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@15107.4 package.scala 96:25:@15108.4]
  assign _T_2509 = _T_2481 ? Mem1D_4_io_output : _T_2508; // @[Mux.scala 31:69:@15171.4]
  assign _T_2478 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@15099.4 package.scala 96:25:@15100.4]
  assign _T_2510 = _T_2478 ? Mem1D_3_io_output : _T_2509; // @[Mux.scala 31:69:@15172.4]
  assign _T_2475 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@15091.4 package.scala 96:25:@15092.4]
  assign _T_2511 = _T_2475 ? Mem1D_2_io_output : _T_2510; // @[Mux.scala 31:69:@15173.4]
  assign _T_2472 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@15083.4 package.scala 96:25:@15084.4]
  assign _T_2512 = _T_2472 ? Mem1D_1_io_output : _T_2511; // @[Mux.scala 31:69:@15174.4]
  assign _T_2469 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@15075.4 package.scala 96:25:@15076.4]
  assign io_rPort_8_output_0 = _T_2469 ? Mem1D_io_output : _T_2512; // @[MemPrimitives.scala 152:13:@15176.4]
  assign io_rPort_7_output_0 = _T_2362 ? Mem1D_io_output : _T_2405; // @[MemPrimitives.scala 152:13:@15032.4]
  assign io_rPort_6_output_0 = _T_2255 ? Mem1D_io_output : _T_2298; // @[MemPrimitives.scala 152:13:@14888.4]
  assign io_rPort_5_output_0 = _T_2148 ? Mem1D_io_output : _T_2191; // @[MemPrimitives.scala 152:13:@14744.4]
  assign io_rPort_4_output_0 = _T_2041 ? Mem1D_io_output : _T_2084; // @[MemPrimitives.scala 152:13:@14600.4]
  assign io_rPort_3_output_0 = _T_1934 ? Mem1D_io_output : _T_1977; // @[MemPrimitives.scala 152:13:@14456.4]
  assign io_rPort_2_output_0 = _T_1827 ? Mem1D_io_output : _T_1870; // @[MemPrimitives.scala 152:13:@14312.4]
  assign io_rPort_1_output_0 = _T_1720 ? Mem1D_io_output : _T_1763; // @[MemPrimitives.scala 152:13:@14168.4]
  assign io_rPort_0_output_0 = _T_1613 ? Mem1D_io_output : _T_1656; // @[MemPrimitives.scala 152:13:@14024.4]
  assign Mem1D_clock = clock; // @[:@12478.4]
  assign Mem1D_reset = reset; // @[:@12479.4]
  assign Mem1D_io_r_ofs_0 = _T_535[9:0]; // @[MemPrimitives.scala 131:28:@12899.4]
  assign Mem1D_io_r_backpressure = _T_535[10]; // @[MemPrimitives.scala 132:32:@12900.4]
  assign Mem1D_io_w_ofs_0 = _T_322[9:0]; // @[MemPrimitives.scala 94:28:@12678.4]
  assign Mem1D_io_w_data_0 = _T_322[41:10]; // @[MemPrimitives.scala 95:29:@12679.4]
  assign Mem1D_io_w_en_0 = _T_322[42]; // @[MemPrimitives.scala 96:27:@12680.4]
  assign Mem1D_1_clock = clock; // @[:@12494.4]
  assign Mem1D_1_reset = reset; // @[:@12495.4]
  assign Mem1D_1_io_r_ofs_0 = _T_627[9:0]; // @[MemPrimitives.scala 131:28:@12988.4]
  assign Mem1D_1_io_r_backpressure = _T_627[10]; // @[MemPrimitives.scala 132:32:@12989.4]
  assign Mem1D_1_io_w_ofs_0 = _T_333[9:0]; // @[MemPrimitives.scala 94:28:@12690.4]
  assign Mem1D_1_io_w_data_0 = _T_333[41:10]; // @[MemPrimitives.scala 95:29:@12691.4]
  assign Mem1D_1_io_w_en_0 = _T_333[42]; // @[MemPrimitives.scala 96:27:@12692.4]
  assign Mem1D_2_clock = clock; // @[:@12510.4]
  assign Mem1D_2_reset = reset; // @[:@12511.4]
  assign Mem1D_2_io_r_ofs_0 = _T_719[9:0]; // @[MemPrimitives.scala 131:28:@13077.4]
  assign Mem1D_2_io_r_backpressure = _T_719[10]; // @[MemPrimitives.scala 132:32:@13078.4]
  assign Mem1D_2_io_w_ofs_0 = _T_344[9:0]; // @[MemPrimitives.scala 94:28:@12702.4]
  assign Mem1D_2_io_w_data_0 = _T_344[41:10]; // @[MemPrimitives.scala 95:29:@12703.4]
  assign Mem1D_2_io_w_en_0 = _T_344[42]; // @[MemPrimitives.scala 96:27:@12704.4]
  assign Mem1D_3_clock = clock; // @[:@12526.4]
  assign Mem1D_3_reset = reset; // @[:@12527.4]
  assign Mem1D_3_io_r_ofs_0 = _T_811[9:0]; // @[MemPrimitives.scala 131:28:@13166.4]
  assign Mem1D_3_io_r_backpressure = _T_811[10]; // @[MemPrimitives.scala 132:32:@13167.4]
  assign Mem1D_3_io_w_ofs_0 = _T_355[9:0]; // @[MemPrimitives.scala 94:28:@12714.4]
  assign Mem1D_3_io_w_data_0 = _T_355[41:10]; // @[MemPrimitives.scala 95:29:@12715.4]
  assign Mem1D_3_io_w_en_0 = _T_355[42]; // @[MemPrimitives.scala 96:27:@12716.4]
  assign Mem1D_4_clock = clock; // @[:@12542.4]
  assign Mem1D_4_reset = reset; // @[:@12543.4]
  assign Mem1D_4_io_r_ofs_0 = _T_903[9:0]; // @[MemPrimitives.scala 131:28:@13255.4]
  assign Mem1D_4_io_r_backpressure = _T_903[10]; // @[MemPrimitives.scala 132:32:@13256.4]
  assign Mem1D_4_io_w_ofs_0 = _T_366[9:0]; // @[MemPrimitives.scala 94:28:@12726.4]
  assign Mem1D_4_io_w_data_0 = _T_366[41:10]; // @[MemPrimitives.scala 95:29:@12727.4]
  assign Mem1D_4_io_w_en_0 = _T_366[42]; // @[MemPrimitives.scala 96:27:@12728.4]
  assign Mem1D_5_clock = clock; // @[:@12558.4]
  assign Mem1D_5_reset = reset; // @[:@12559.4]
  assign Mem1D_5_io_r_ofs_0 = _T_995[9:0]; // @[MemPrimitives.scala 131:28:@13344.4]
  assign Mem1D_5_io_r_backpressure = _T_995[10]; // @[MemPrimitives.scala 132:32:@13345.4]
  assign Mem1D_5_io_w_ofs_0 = _T_377[9:0]; // @[MemPrimitives.scala 94:28:@12738.4]
  assign Mem1D_5_io_w_data_0 = _T_377[41:10]; // @[MemPrimitives.scala 95:29:@12739.4]
  assign Mem1D_5_io_w_en_0 = _T_377[42]; // @[MemPrimitives.scala 96:27:@12740.4]
  assign Mem1D_6_clock = clock; // @[:@12574.4]
  assign Mem1D_6_reset = reset; // @[:@12575.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1087[9:0]; // @[MemPrimitives.scala 131:28:@13433.4]
  assign Mem1D_6_io_r_backpressure = _T_1087[10]; // @[MemPrimitives.scala 132:32:@13434.4]
  assign Mem1D_6_io_w_ofs_0 = _T_388[9:0]; // @[MemPrimitives.scala 94:28:@12750.4]
  assign Mem1D_6_io_w_data_0 = _T_388[41:10]; // @[MemPrimitives.scala 95:29:@12751.4]
  assign Mem1D_6_io_w_en_0 = _T_388[42]; // @[MemPrimitives.scala 96:27:@12752.4]
  assign Mem1D_7_clock = clock; // @[:@12590.4]
  assign Mem1D_7_reset = reset; // @[:@12591.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1179[9:0]; // @[MemPrimitives.scala 131:28:@13522.4]
  assign Mem1D_7_io_r_backpressure = _T_1179[10]; // @[MemPrimitives.scala 132:32:@13523.4]
  assign Mem1D_7_io_w_ofs_0 = _T_399[9:0]; // @[MemPrimitives.scala 94:28:@12762.4]
  assign Mem1D_7_io_w_data_0 = _T_399[41:10]; // @[MemPrimitives.scala 95:29:@12763.4]
  assign Mem1D_7_io_w_en_0 = _T_399[42]; // @[MemPrimitives.scala 96:27:@12764.4]
  assign Mem1D_8_clock = clock; // @[:@12606.4]
  assign Mem1D_8_reset = reset; // @[:@12607.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1271[9:0]; // @[MemPrimitives.scala 131:28:@13611.4]
  assign Mem1D_8_io_r_backpressure = _T_1271[10]; // @[MemPrimitives.scala 132:32:@13612.4]
  assign Mem1D_8_io_w_ofs_0 = _T_410[9:0]; // @[MemPrimitives.scala 94:28:@12774.4]
  assign Mem1D_8_io_w_data_0 = _T_410[41:10]; // @[MemPrimitives.scala 95:29:@12775.4]
  assign Mem1D_8_io_w_en_0 = _T_410[42]; // @[MemPrimitives.scala 96:27:@12776.4]
  assign Mem1D_9_clock = clock; // @[:@12622.4]
  assign Mem1D_9_reset = reset; // @[:@12623.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1363[9:0]; // @[MemPrimitives.scala 131:28:@13700.4]
  assign Mem1D_9_io_r_backpressure = _T_1363[10]; // @[MemPrimitives.scala 132:32:@13701.4]
  assign Mem1D_9_io_w_ofs_0 = _T_421[9:0]; // @[MemPrimitives.scala 94:28:@12786.4]
  assign Mem1D_9_io_w_data_0 = _T_421[41:10]; // @[MemPrimitives.scala 95:29:@12787.4]
  assign Mem1D_9_io_w_en_0 = _T_421[42]; // @[MemPrimitives.scala 96:27:@12788.4]
  assign Mem1D_10_clock = clock; // @[:@12638.4]
  assign Mem1D_10_reset = reset; // @[:@12639.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1455[9:0]; // @[MemPrimitives.scala 131:28:@13789.4]
  assign Mem1D_10_io_r_backpressure = _T_1455[10]; // @[MemPrimitives.scala 132:32:@13790.4]
  assign Mem1D_10_io_w_ofs_0 = _T_432[9:0]; // @[MemPrimitives.scala 94:28:@12798.4]
  assign Mem1D_10_io_w_data_0 = _T_432[41:10]; // @[MemPrimitives.scala 95:29:@12799.4]
  assign Mem1D_10_io_w_en_0 = _T_432[42]; // @[MemPrimitives.scala 96:27:@12800.4]
  assign Mem1D_11_clock = clock; // @[:@12654.4]
  assign Mem1D_11_reset = reset; // @[:@12655.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1547[9:0]; // @[MemPrimitives.scala 131:28:@13878.4]
  assign Mem1D_11_io_r_backpressure = _T_1547[10]; // @[MemPrimitives.scala 132:32:@13879.4]
  assign Mem1D_11_io_w_ofs_0 = _T_443[9:0]; // @[MemPrimitives.scala 94:28:@12810.4]
  assign Mem1D_11_io_w_data_0 = _T_443[41:10]; // @[MemPrimitives.scala 95:29:@12811.4]
  assign Mem1D_11_io_w_en_0 = _T_443[42]; // @[MemPrimitives.scala 96:27:@12812.4]
  assign StickySelects_clock = clock; // @[:@12850.4]
  assign StickySelects_reset = reset; // @[:@12851.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_451; // @[MemPrimitives.scala 125:64:@12852.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_457; // @[MemPrimitives.scala 125:64:@12853.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_463; // @[MemPrimitives.scala 125:64:@12854.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_469; // @[MemPrimitives.scala 125:64:@12855.4]
  assign StickySelects_io_ins_4 = io_rPort_4_en_0 & _T_475; // @[MemPrimitives.scala 125:64:@12856.4]
  assign StickySelects_io_ins_5 = io_rPort_5_en_0 & _T_481; // @[MemPrimitives.scala 125:64:@12857.4]
  assign StickySelects_io_ins_6 = io_rPort_6_en_0 & _T_487; // @[MemPrimitives.scala 125:64:@12858.4]
  assign StickySelects_io_ins_7 = io_rPort_7_en_0 & _T_493; // @[MemPrimitives.scala 125:64:@12859.4]
  assign StickySelects_io_ins_8 = io_rPort_8_en_0 & _T_499; // @[MemPrimitives.scala 125:64:@12860.4]
  assign StickySelects_1_clock = clock; // @[:@12939.4]
  assign StickySelects_1_reset = reset; // @[:@12940.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_543; // @[MemPrimitives.scala 125:64:@12941.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_549; // @[MemPrimitives.scala 125:64:@12942.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_555; // @[MemPrimitives.scala 125:64:@12943.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_561; // @[MemPrimitives.scala 125:64:@12944.4]
  assign StickySelects_1_io_ins_4 = io_rPort_4_en_0 & _T_567; // @[MemPrimitives.scala 125:64:@12945.4]
  assign StickySelects_1_io_ins_5 = io_rPort_5_en_0 & _T_573; // @[MemPrimitives.scala 125:64:@12946.4]
  assign StickySelects_1_io_ins_6 = io_rPort_6_en_0 & _T_579; // @[MemPrimitives.scala 125:64:@12947.4]
  assign StickySelects_1_io_ins_7 = io_rPort_7_en_0 & _T_585; // @[MemPrimitives.scala 125:64:@12948.4]
  assign StickySelects_1_io_ins_8 = io_rPort_8_en_0 & _T_591; // @[MemPrimitives.scala 125:64:@12949.4]
  assign StickySelects_2_clock = clock; // @[:@13028.4]
  assign StickySelects_2_reset = reset; // @[:@13029.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@13030.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@13031.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@13032.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@13033.4]
  assign StickySelects_2_io_ins_4 = io_rPort_4_en_0 & _T_659; // @[MemPrimitives.scala 125:64:@13034.4]
  assign StickySelects_2_io_ins_5 = io_rPort_5_en_0 & _T_665; // @[MemPrimitives.scala 125:64:@13035.4]
  assign StickySelects_2_io_ins_6 = io_rPort_6_en_0 & _T_671; // @[MemPrimitives.scala 125:64:@13036.4]
  assign StickySelects_2_io_ins_7 = io_rPort_7_en_0 & _T_677; // @[MemPrimitives.scala 125:64:@13037.4]
  assign StickySelects_2_io_ins_8 = io_rPort_8_en_0 & _T_683; // @[MemPrimitives.scala 125:64:@13038.4]
  assign StickySelects_3_clock = clock; // @[:@13117.4]
  assign StickySelects_3_reset = reset; // @[:@13118.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@13119.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@13120.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@13121.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_745; // @[MemPrimitives.scala 125:64:@13122.4]
  assign StickySelects_3_io_ins_4 = io_rPort_4_en_0 & _T_751; // @[MemPrimitives.scala 125:64:@13123.4]
  assign StickySelects_3_io_ins_5 = io_rPort_5_en_0 & _T_757; // @[MemPrimitives.scala 125:64:@13124.4]
  assign StickySelects_3_io_ins_6 = io_rPort_6_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@13125.4]
  assign StickySelects_3_io_ins_7 = io_rPort_7_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@13126.4]
  assign StickySelects_3_io_ins_8 = io_rPort_8_en_0 & _T_775; // @[MemPrimitives.scala 125:64:@13127.4]
  assign StickySelects_4_clock = clock; // @[:@13206.4]
  assign StickySelects_4_reset = reset; // @[:@13207.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_819; // @[MemPrimitives.scala 125:64:@13208.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_825; // @[MemPrimitives.scala 125:64:@13209.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_831; // @[MemPrimitives.scala 125:64:@13210.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_837; // @[MemPrimitives.scala 125:64:@13211.4]
  assign StickySelects_4_io_ins_4 = io_rPort_4_en_0 & _T_843; // @[MemPrimitives.scala 125:64:@13212.4]
  assign StickySelects_4_io_ins_5 = io_rPort_5_en_0 & _T_849; // @[MemPrimitives.scala 125:64:@13213.4]
  assign StickySelects_4_io_ins_6 = io_rPort_6_en_0 & _T_855; // @[MemPrimitives.scala 125:64:@13214.4]
  assign StickySelects_4_io_ins_7 = io_rPort_7_en_0 & _T_861; // @[MemPrimitives.scala 125:64:@13215.4]
  assign StickySelects_4_io_ins_8 = io_rPort_8_en_0 & _T_867; // @[MemPrimitives.scala 125:64:@13216.4]
  assign StickySelects_5_clock = clock; // @[:@13295.4]
  assign StickySelects_5_reset = reset; // @[:@13296.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_911; // @[MemPrimitives.scala 125:64:@13297.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_917; // @[MemPrimitives.scala 125:64:@13298.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_923; // @[MemPrimitives.scala 125:64:@13299.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_929; // @[MemPrimitives.scala 125:64:@13300.4]
  assign StickySelects_5_io_ins_4 = io_rPort_4_en_0 & _T_935; // @[MemPrimitives.scala 125:64:@13301.4]
  assign StickySelects_5_io_ins_5 = io_rPort_5_en_0 & _T_941; // @[MemPrimitives.scala 125:64:@13302.4]
  assign StickySelects_5_io_ins_6 = io_rPort_6_en_0 & _T_947; // @[MemPrimitives.scala 125:64:@13303.4]
  assign StickySelects_5_io_ins_7 = io_rPort_7_en_0 & _T_953; // @[MemPrimitives.scala 125:64:@13304.4]
  assign StickySelects_5_io_ins_8 = io_rPort_8_en_0 & _T_959; // @[MemPrimitives.scala 125:64:@13305.4]
  assign StickySelects_6_clock = clock; // @[:@13384.4]
  assign StickySelects_6_reset = reset; // @[:@13385.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1003; // @[MemPrimitives.scala 125:64:@13386.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1009; // @[MemPrimitives.scala 125:64:@13387.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_1015; // @[MemPrimitives.scala 125:64:@13388.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_1021; // @[MemPrimitives.scala 125:64:@13389.4]
  assign StickySelects_6_io_ins_4 = io_rPort_4_en_0 & _T_1027; // @[MemPrimitives.scala 125:64:@13390.4]
  assign StickySelects_6_io_ins_5 = io_rPort_5_en_0 & _T_1033; // @[MemPrimitives.scala 125:64:@13391.4]
  assign StickySelects_6_io_ins_6 = io_rPort_6_en_0 & _T_1039; // @[MemPrimitives.scala 125:64:@13392.4]
  assign StickySelects_6_io_ins_7 = io_rPort_7_en_0 & _T_1045; // @[MemPrimitives.scala 125:64:@13393.4]
  assign StickySelects_6_io_ins_8 = io_rPort_8_en_0 & _T_1051; // @[MemPrimitives.scala 125:64:@13394.4]
  assign StickySelects_7_clock = clock; // @[:@13473.4]
  assign StickySelects_7_reset = reset; // @[:@13474.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1095; // @[MemPrimitives.scala 125:64:@13475.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1101; // @[MemPrimitives.scala 125:64:@13476.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1107; // @[MemPrimitives.scala 125:64:@13477.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1113; // @[MemPrimitives.scala 125:64:@13478.4]
  assign StickySelects_7_io_ins_4 = io_rPort_4_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13479.4]
  assign StickySelects_7_io_ins_5 = io_rPort_5_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13480.4]
  assign StickySelects_7_io_ins_6 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13481.4]
  assign StickySelects_7_io_ins_7 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13482.4]
  assign StickySelects_7_io_ins_8 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13483.4]
  assign StickySelects_8_clock = clock; // @[:@13562.4]
  assign StickySelects_8_reset = reset; // @[:@13563.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13564.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13565.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13566.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13567.4]
  assign StickySelects_8_io_ins_4 = io_rPort_4_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13568.4]
  assign StickySelects_8_io_ins_5 = io_rPort_5_en_0 & _T_1217; // @[MemPrimitives.scala 125:64:@13569.4]
  assign StickySelects_8_io_ins_6 = io_rPort_6_en_0 & _T_1223; // @[MemPrimitives.scala 125:64:@13570.4]
  assign StickySelects_8_io_ins_7 = io_rPort_7_en_0 & _T_1229; // @[MemPrimitives.scala 125:64:@13571.4]
  assign StickySelects_8_io_ins_8 = io_rPort_8_en_0 & _T_1235; // @[MemPrimitives.scala 125:64:@13572.4]
  assign StickySelects_9_clock = clock; // @[:@13651.4]
  assign StickySelects_9_reset = reset; // @[:@13652.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1279; // @[MemPrimitives.scala 125:64:@13653.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1285; // @[MemPrimitives.scala 125:64:@13654.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1291; // @[MemPrimitives.scala 125:64:@13655.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1297; // @[MemPrimitives.scala 125:64:@13656.4]
  assign StickySelects_9_io_ins_4 = io_rPort_4_en_0 & _T_1303; // @[MemPrimitives.scala 125:64:@13657.4]
  assign StickySelects_9_io_ins_5 = io_rPort_5_en_0 & _T_1309; // @[MemPrimitives.scala 125:64:@13658.4]
  assign StickySelects_9_io_ins_6 = io_rPort_6_en_0 & _T_1315; // @[MemPrimitives.scala 125:64:@13659.4]
  assign StickySelects_9_io_ins_7 = io_rPort_7_en_0 & _T_1321; // @[MemPrimitives.scala 125:64:@13660.4]
  assign StickySelects_9_io_ins_8 = io_rPort_8_en_0 & _T_1327; // @[MemPrimitives.scala 125:64:@13661.4]
  assign StickySelects_10_clock = clock; // @[:@13740.4]
  assign StickySelects_10_reset = reset; // @[:@13741.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1371; // @[MemPrimitives.scala 125:64:@13742.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_1377; // @[MemPrimitives.scala 125:64:@13743.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_1383; // @[MemPrimitives.scala 125:64:@13744.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_1389; // @[MemPrimitives.scala 125:64:@13745.4]
  assign StickySelects_10_io_ins_4 = io_rPort_4_en_0 & _T_1395; // @[MemPrimitives.scala 125:64:@13746.4]
  assign StickySelects_10_io_ins_5 = io_rPort_5_en_0 & _T_1401; // @[MemPrimitives.scala 125:64:@13747.4]
  assign StickySelects_10_io_ins_6 = io_rPort_6_en_0 & _T_1407; // @[MemPrimitives.scala 125:64:@13748.4]
  assign StickySelects_10_io_ins_7 = io_rPort_7_en_0 & _T_1413; // @[MemPrimitives.scala 125:64:@13749.4]
  assign StickySelects_10_io_ins_8 = io_rPort_8_en_0 & _T_1419; // @[MemPrimitives.scala 125:64:@13750.4]
  assign StickySelects_11_clock = clock; // @[:@13829.4]
  assign StickySelects_11_reset = reset; // @[:@13830.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1463; // @[MemPrimitives.scala 125:64:@13831.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1469; // @[MemPrimitives.scala 125:64:@13832.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1475; // @[MemPrimitives.scala 125:64:@13833.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1481; // @[MemPrimitives.scala 125:64:@13834.4]
  assign StickySelects_11_io_ins_4 = io_rPort_4_en_0 & _T_1487; // @[MemPrimitives.scala 125:64:@13835.4]
  assign StickySelects_11_io_ins_5 = io_rPort_5_en_0 & _T_1493; // @[MemPrimitives.scala 125:64:@13836.4]
  assign StickySelects_11_io_ins_6 = io_rPort_6_en_0 & _T_1499; // @[MemPrimitives.scala 125:64:@13837.4]
  assign StickySelects_11_io_ins_7 = io_rPort_7_en_0 & _T_1505; // @[MemPrimitives.scala 125:64:@13838.4]
  assign StickySelects_11_io_ins_8 = io_rPort_8_en_0 & _T_1511; // @[MemPrimitives.scala 125:64:@13839.4]
  assign RetimeWrapper_clock = clock; // @[:@13919.4]
  assign RetimeWrapper_reset = reset; // @[:@13920.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13922.4]
  assign RetimeWrapper_io_in = _T_451 & io_rPort_0_en_0; // @[package.scala 94:16:@13921.4]
  assign RetimeWrapper_1_clock = clock; // @[:@13927.4]
  assign RetimeWrapper_1_reset = reset; // @[:@13928.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13930.4]
  assign RetimeWrapper_1_io_in = _T_543 & io_rPort_0_en_0; // @[package.scala 94:16:@13929.4]
  assign RetimeWrapper_2_clock = clock; // @[:@13935.4]
  assign RetimeWrapper_2_reset = reset; // @[:@13936.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13938.4]
  assign RetimeWrapper_2_io_in = _T_635 & io_rPort_0_en_0; // @[package.scala 94:16:@13937.4]
  assign RetimeWrapper_3_clock = clock; // @[:@13943.4]
  assign RetimeWrapper_3_reset = reset; // @[:@13944.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13946.4]
  assign RetimeWrapper_3_io_in = _T_727 & io_rPort_0_en_0; // @[package.scala 94:16:@13945.4]
  assign RetimeWrapper_4_clock = clock; // @[:@13951.4]
  assign RetimeWrapper_4_reset = reset; // @[:@13952.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13954.4]
  assign RetimeWrapper_4_io_in = _T_819 & io_rPort_0_en_0; // @[package.scala 94:16:@13953.4]
  assign RetimeWrapper_5_clock = clock; // @[:@13959.4]
  assign RetimeWrapper_5_reset = reset; // @[:@13960.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13962.4]
  assign RetimeWrapper_5_io_in = _T_911 & io_rPort_0_en_0; // @[package.scala 94:16:@13961.4]
  assign RetimeWrapper_6_clock = clock; // @[:@13967.4]
  assign RetimeWrapper_6_reset = reset; // @[:@13968.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13970.4]
  assign RetimeWrapper_6_io_in = _T_1003 & io_rPort_0_en_0; // @[package.scala 94:16:@13969.4]
  assign RetimeWrapper_7_clock = clock; // @[:@13975.4]
  assign RetimeWrapper_7_reset = reset; // @[:@13976.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13978.4]
  assign RetimeWrapper_7_io_in = _T_1095 & io_rPort_0_en_0; // @[package.scala 94:16:@13977.4]
  assign RetimeWrapper_8_clock = clock; // @[:@13983.4]
  assign RetimeWrapper_8_reset = reset; // @[:@13984.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13986.4]
  assign RetimeWrapper_8_io_in = _T_1187 & io_rPort_0_en_0; // @[package.scala 94:16:@13985.4]
  assign RetimeWrapper_9_clock = clock; // @[:@13991.4]
  assign RetimeWrapper_9_reset = reset; // @[:@13992.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13994.4]
  assign RetimeWrapper_9_io_in = _T_1279 & io_rPort_0_en_0; // @[package.scala 94:16:@13993.4]
  assign RetimeWrapper_10_clock = clock; // @[:@13999.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14000.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14002.4]
  assign RetimeWrapper_10_io_in = _T_1371 & io_rPort_0_en_0; // @[package.scala 94:16:@14001.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14007.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14008.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14010.4]
  assign RetimeWrapper_11_io_in = _T_1463 & io_rPort_0_en_0; // @[package.scala 94:16:@14009.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14063.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14064.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14066.4]
  assign RetimeWrapper_12_io_in = _T_457 & io_rPort_1_en_0; // @[package.scala 94:16:@14065.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14071.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14072.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14074.4]
  assign RetimeWrapper_13_io_in = _T_549 & io_rPort_1_en_0; // @[package.scala 94:16:@14073.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14079.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14080.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14082.4]
  assign RetimeWrapper_14_io_in = _T_641 & io_rPort_1_en_0; // @[package.scala 94:16:@14081.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14087.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14088.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14090.4]
  assign RetimeWrapper_15_io_in = _T_733 & io_rPort_1_en_0; // @[package.scala 94:16:@14089.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14095.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14096.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14098.4]
  assign RetimeWrapper_16_io_in = _T_825 & io_rPort_1_en_0; // @[package.scala 94:16:@14097.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14103.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14104.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14106.4]
  assign RetimeWrapper_17_io_in = _T_917 & io_rPort_1_en_0; // @[package.scala 94:16:@14105.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14111.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14112.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14114.4]
  assign RetimeWrapper_18_io_in = _T_1009 & io_rPort_1_en_0; // @[package.scala 94:16:@14113.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14119.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14120.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14122.4]
  assign RetimeWrapper_19_io_in = _T_1101 & io_rPort_1_en_0; // @[package.scala 94:16:@14121.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14127.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14128.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14130.4]
  assign RetimeWrapper_20_io_in = _T_1193 & io_rPort_1_en_0; // @[package.scala 94:16:@14129.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14135.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14136.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14138.4]
  assign RetimeWrapper_21_io_in = _T_1285 & io_rPort_1_en_0; // @[package.scala 94:16:@14137.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14143.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14144.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14146.4]
  assign RetimeWrapper_22_io_in = _T_1377 & io_rPort_1_en_0; // @[package.scala 94:16:@14145.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14151.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14152.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14154.4]
  assign RetimeWrapper_23_io_in = _T_1469 & io_rPort_1_en_0; // @[package.scala 94:16:@14153.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14207.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14208.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14210.4]
  assign RetimeWrapper_24_io_in = _T_463 & io_rPort_2_en_0; // @[package.scala 94:16:@14209.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14215.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14216.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14218.4]
  assign RetimeWrapper_25_io_in = _T_555 & io_rPort_2_en_0; // @[package.scala 94:16:@14217.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14223.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14224.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14226.4]
  assign RetimeWrapper_26_io_in = _T_647 & io_rPort_2_en_0; // @[package.scala 94:16:@14225.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14231.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14232.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14234.4]
  assign RetimeWrapper_27_io_in = _T_739 & io_rPort_2_en_0; // @[package.scala 94:16:@14233.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14239.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14240.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14242.4]
  assign RetimeWrapper_28_io_in = _T_831 & io_rPort_2_en_0; // @[package.scala 94:16:@14241.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14247.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14248.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14250.4]
  assign RetimeWrapper_29_io_in = _T_923 & io_rPort_2_en_0; // @[package.scala 94:16:@14249.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14255.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14256.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14258.4]
  assign RetimeWrapper_30_io_in = _T_1015 & io_rPort_2_en_0; // @[package.scala 94:16:@14257.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14263.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14264.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14266.4]
  assign RetimeWrapper_31_io_in = _T_1107 & io_rPort_2_en_0; // @[package.scala 94:16:@14265.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14271.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14272.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14274.4]
  assign RetimeWrapper_32_io_in = _T_1199 & io_rPort_2_en_0; // @[package.scala 94:16:@14273.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14279.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14280.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14282.4]
  assign RetimeWrapper_33_io_in = _T_1291 & io_rPort_2_en_0; // @[package.scala 94:16:@14281.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14287.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14288.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14290.4]
  assign RetimeWrapper_34_io_in = _T_1383 & io_rPort_2_en_0; // @[package.scala 94:16:@14289.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14295.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14296.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14298.4]
  assign RetimeWrapper_35_io_in = _T_1475 & io_rPort_2_en_0; // @[package.scala 94:16:@14297.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14351.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14352.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14354.4]
  assign RetimeWrapper_36_io_in = _T_469 & io_rPort_3_en_0; // @[package.scala 94:16:@14353.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14359.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14360.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14362.4]
  assign RetimeWrapper_37_io_in = _T_561 & io_rPort_3_en_0; // @[package.scala 94:16:@14361.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14367.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14368.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14370.4]
  assign RetimeWrapper_38_io_in = _T_653 & io_rPort_3_en_0; // @[package.scala 94:16:@14369.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14375.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14376.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14378.4]
  assign RetimeWrapper_39_io_in = _T_745 & io_rPort_3_en_0; // @[package.scala 94:16:@14377.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14383.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14384.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14386.4]
  assign RetimeWrapper_40_io_in = _T_837 & io_rPort_3_en_0; // @[package.scala 94:16:@14385.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14391.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14392.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14394.4]
  assign RetimeWrapper_41_io_in = _T_929 & io_rPort_3_en_0; // @[package.scala 94:16:@14393.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14399.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14400.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14402.4]
  assign RetimeWrapper_42_io_in = _T_1021 & io_rPort_3_en_0; // @[package.scala 94:16:@14401.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14407.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14408.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14410.4]
  assign RetimeWrapper_43_io_in = _T_1113 & io_rPort_3_en_0; // @[package.scala 94:16:@14409.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14415.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14416.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14418.4]
  assign RetimeWrapper_44_io_in = _T_1205 & io_rPort_3_en_0; // @[package.scala 94:16:@14417.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14423.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14424.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14426.4]
  assign RetimeWrapper_45_io_in = _T_1297 & io_rPort_3_en_0; // @[package.scala 94:16:@14425.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14431.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14432.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14434.4]
  assign RetimeWrapper_46_io_in = _T_1389 & io_rPort_3_en_0; // @[package.scala 94:16:@14433.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14439.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14440.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14442.4]
  assign RetimeWrapper_47_io_in = _T_1481 & io_rPort_3_en_0; // @[package.scala 94:16:@14441.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14495.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14496.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14498.4]
  assign RetimeWrapper_48_io_in = _T_475 & io_rPort_4_en_0; // @[package.scala 94:16:@14497.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14503.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14504.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14506.4]
  assign RetimeWrapper_49_io_in = _T_567 & io_rPort_4_en_0; // @[package.scala 94:16:@14505.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14511.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14512.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14514.4]
  assign RetimeWrapper_50_io_in = _T_659 & io_rPort_4_en_0; // @[package.scala 94:16:@14513.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14519.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14520.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14522.4]
  assign RetimeWrapper_51_io_in = _T_751 & io_rPort_4_en_0; // @[package.scala 94:16:@14521.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14527.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14528.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14530.4]
  assign RetimeWrapper_52_io_in = _T_843 & io_rPort_4_en_0; // @[package.scala 94:16:@14529.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14535.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14536.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14538.4]
  assign RetimeWrapper_53_io_in = _T_935 & io_rPort_4_en_0; // @[package.scala 94:16:@14537.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14543.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14544.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14546.4]
  assign RetimeWrapper_54_io_in = _T_1027 & io_rPort_4_en_0; // @[package.scala 94:16:@14545.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14551.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14552.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14554.4]
  assign RetimeWrapper_55_io_in = _T_1119 & io_rPort_4_en_0; // @[package.scala 94:16:@14553.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14559.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14560.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14562.4]
  assign RetimeWrapper_56_io_in = _T_1211 & io_rPort_4_en_0; // @[package.scala 94:16:@14561.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14567.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14568.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14570.4]
  assign RetimeWrapper_57_io_in = _T_1303 & io_rPort_4_en_0; // @[package.scala 94:16:@14569.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14575.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14576.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14578.4]
  assign RetimeWrapper_58_io_in = _T_1395 & io_rPort_4_en_0; // @[package.scala 94:16:@14577.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14583.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14584.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14586.4]
  assign RetimeWrapper_59_io_in = _T_1487 & io_rPort_4_en_0; // @[package.scala 94:16:@14585.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14639.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14640.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14642.4]
  assign RetimeWrapper_60_io_in = _T_481 & io_rPort_5_en_0; // @[package.scala 94:16:@14641.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14647.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14648.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14650.4]
  assign RetimeWrapper_61_io_in = _T_573 & io_rPort_5_en_0; // @[package.scala 94:16:@14649.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14655.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14656.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14658.4]
  assign RetimeWrapper_62_io_in = _T_665 & io_rPort_5_en_0; // @[package.scala 94:16:@14657.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14663.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14664.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14666.4]
  assign RetimeWrapper_63_io_in = _T_757 & io_rPort_5_en_0; // @[package.scala 94:16:@14665.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14671.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14672.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14674.4]
  assign RetimeWrapper_64_io_in = _T_849 & io_rPort_5_en_0; // @[package.scala 94:16:@14673.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14679.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14680.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14682.4]
  assign RetimeWrapper_65_io_in = _T_941 & io_rPort_5_en_0; // @[package.scala 94:16:@14681.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14687.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14688.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14690.4]
  assign RetimeWrapper_66_io_in = _T_1033 & io_rPort_5_en_0; // @[package.scala 94:16:@14689.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14695.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14696.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14698.4]
  assign RetimeWrapper_67_io_in = _T_1125 & io_rPort_5_en_0; // @[package.scala 94:16:@14697.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14703.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14704.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14706.4]
  assign RetimeWrapper_68_io_in = _T_1217 & io_rPort_5_en_0; // @[package.scala 94:16:@14705.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14711.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14712.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14714.4]
  assign RetimeWrapper_69_io_in = _T_1309 & io_rPort_5_en_0; // @[package.scala 94:16:@14713.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14719.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14720.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14722.4]
  assign RetimeWrapper_70_io_in = _T_1401 & io_rPort_5_en_0; // @[package.scala 94:16:@14721.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14727.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14728.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14730.4]
  assign RetimeWrapper_71_io_in = _T_1493 & io_rPort_5_en_0; // @[package.scala 94:16:@14729.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14783.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14784.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14786.4]
  assign RetimeWrapper_72_io_in = _T_487 & io_rPort_6_en_0; // @[package.scala 94:16:@14785.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14791.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14792.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14794.4]
  assign RetimeWrapper_73_io_in = _T_579 & io_rPort_6_en_0; // @[package.scala 94:16:@14793.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14799.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14800.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14802.4]
  assign RetimeWrapper_74_io_in = _T_671 & io_rPort_6_en_0; // @[package.scala 94:16:@14801.4]
  assign RetimeWrapper_75_clock = clock; // @[:@14807.4]
  assign RetimeWrapper_75_reset = reset; // @[:@14808.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14810.4]
  assign RetimeWrapper_75_io_in = _T_763 & io_rPort_6_en_0; // @[package.scala 94:16:@14809.4]
  assign RetimeWrapper_76_clock = clock; // @[:@14815.4]
  assign RetimeWrapper_76_reset = reset; // @[:@14816.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14818.4]
  assign RetimeWrapper_76_io_in = _T_855 & io_rPort_6_en_0; // @[package.scala 94:16:@14817.4]
  assign RetimeWrapper_77_clock = clock; // @[:@14823.4]
  assign RetimeWrapper_77_reset = reset; // @[:@14824.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14826.4]
  assign RetimeWrapper_77_io_in = _T_947 & io_rPort_6_en_0; // @[package.scala 94:16:@14825.4]
  assign RetimeWrapper_78_clock = clock; // @[:@14831.4]
  assign RetimeWrapper_78_reset = reset; // @[:@14832.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14834.4]
  assign RetimeWrapper_78_io_in = _T_1039 & io_rPort_6_en_0; // @[package.scala 94:16:@14833.4]
  assign RetimeWrapper_79_clock = clock; // @[:@14839.4]
  assign RetimeWrapper_79_reset = reset; // @[:@14840.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14842.4]
  assign RetimeWrapper_79_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@14841.4]
  assign RetimeWrapper_80_clock = clock; // @[:@14847.4]
  assign RetimeWrapper_80_reset = reset; // @[:@14848.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14850.4]
  assign RetimeWrapper_80_io_in = _T_1223 & io_rPort_6_en_0; // @[package.scala 94:16:@14849.4]
  assign RetimeWrapper_81_clock = clock; // @[:@14855.4]
  assign RetimeWrapper_81_reset = reset; // @[:@14856.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14858.4]
  assign RetimeWrapper_81_io_in = _T_1315 & io_rPort_6_en_0; // @[package.scala 94:16:@14857.4]
  assign RetimeWrapper_82_clock = clock; // @[:@14863.4]
  assign RetimeWrapper_82_reset = reset; // @[:@14864.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14866.4]
  assign RetimeWrapper_82_io_in = _T_1407 & io_rPort_6_en_0; // @[package.scala 94:16:@14865.4]
  assign RetimeWrapper_83_clock = clock; // @[:@14871.4]
  assign RetimeWrapper_83_reset = reset; // @[:@14872.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14874.4]
  assign RetimeWrapper_83_io_in = _T_1499 & io_rPort_6_en_0; // @[package.scala 94:16:@14873.4]
  assign RetimeWrapper_84_clock = clock; // @[:@14927.4]
  assign RetimeWrapper_84_reset = reset; // @[:@14928.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14930.4]
  assign RetimeWrapper_84_io_in = _T_493 & io_rPort_7_en_0; // @[package.scala 94:16:@14929.4]
  assign RetimeWrapper_85_clock = clock; // @[:@14935.4]
  assign RetimeWrapper_85_reset = reset; // @[:@14936.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14938.4]
  assign RetimeWrapper_85_io_in = _T_585 & io_rPort_7_en_0; // @[package.scala 94:16:@14937.4]
  assign RetimeWrapper_86_clock = clock; // @[:@14943.4]
  assign RetimeWrapper_86_reset = reset; // @[:@14944.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14946.4]
  assign RetimeWrapper_86_io_in = _T_677 & io_rPort_7_en_0; // @[package.scala 94:16:@14945.4]
  assign RetimeWrapper_87_clock = clock; // @[:@14951.4]
  assign RetimeWrapper_87_reset = reset; // @[:@14952.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14954.4]
  assign RetimeWrapper_87_io_in = _T_769 & io_rPort_7_en_0; // @[package.scala 94:16:@14953.4]
  assign RetimeWrapper_88_clock = clock; // @[:@14959.4]
  assign RetimeWrapper_88_reset = reset; // @[:@14960.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14962.4]
  assign RetimeWrapper_88_io_in = _T_861 & io_rPort_7_en_0; // @[package.scala 94:16:@14961.4]
  assign RetimeWrapper_89_clock = clock; // @[:@14967.4]
  assign RetimeWrapper_89_reset = reset; // @[:@14968.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14970.4]
  assign RetimeWrapper_89_io_in = _T_953 & io_rPort_7_en_0; // @[package.scala 94:16:@14969.4]
  assign RetimeWrapper_90_clock = clock; // @[:@14975.4]
  assign RetimeWrapper_90_reset = reset; // @[:@14976.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14978.4]
  assign RetimeWrapper_90_io_in = _T_1045 & io_rPort_7_en_0; // @[package.scala 94:16:@14977.4]
  assign RetimeWrapper_91_clock = clock; // @[:@14983.4]
  assign RetimeWrapper_91_reset = reset; // @[:@14984.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14986.4]
  assign RetimeWrapper_91_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@14985.4]
  assign RetimeWrapper_92_clock = clock; // @[:@14991.4]
  assign RetimeWrapper_92_reset = reset; // @[:@14992.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14994.4]
  assign RetimeWrapper_92_io_in = _T_1229 & io_rPort_7_en_0; // @[package.scala 94:16:@14993.4]
  assign RetimeWrapper_93_clock = clock; // @[:@14999.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15000.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15002.4]
  assign RetimeWrapper_93_io_in = _T_1321 & io_rPort_7_en_0; // @[package.scala 94:16:@15001.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15007.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15008.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15010.4]
  assign RetimeWrapper_94_io_in = _T_1413 & io_rPort_7_en_0; // @[package.scala 94:16:@15009.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15015.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15016.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15018.4]
  assign RetimeWrapper_95_io_in = _T_1505 & io_rPort_7_en_0; // @[package.scala 94:16:@15017.4]
  assign RetimeWrapper_96_clock = clock; // @[:@15071.4]
  assign RetimeWrapper_96_reset = reset; // @[:@15072.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15074.4]
  assign RetimeWrapper_96_io_in = _T_499 & io_rPort_8_en_0; // @[package.scala 94:16:@15073.4]
  assign RetimeWrapper_97_clock = clock; // @[:@15079.4]
  assign RetimeWrapper_97_reset = reset; // @[:@15080.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15082.4]
  assign RetimeWrapper_97_io_in = _T_591 & io_rPort_8_en_0; // @[package.scala 94:16:@15081.4]
  assign RetimeWrapper_98_clock = clock; // @[:@15087.4]
  assign RetimeWrapper_98_reset = reset; // @[:@15088.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15090.4]
  assign RetimeWrapper_98_io_in = _T_683 & io_rPort_8_en_0; // @[package.scala 94:16:@15089.4]
  assign RetimeWrapper_99_clock = clock; // @[:@15095.4]
  assign RetimeWrapper_99_reset = reset; // @[:@15096.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15098.4]
  assign RetimeWrapper_99_io_in = _T_775 & io_rPort_8_en_0; // @[package.scala 94:16:@15097.4]
  assign RetimeWrapper_100_clock = clock; // @[:@15103.4]
  assign RetimeWrapper_100_reset = reset; // @[:@15104.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15106.4]
  assign RetimeWrapper_100_io_in = _T_867 & io_rPort_8_en_0; // @[package.scala 94:16:@15105.4]
  assign RetimeWrapper_101_clock = clock; // @[:@15111.4]
  assign RetimeWrapper_101_reset = reset; // @[:@15112.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15114.4]
  assign RetimeWrapper_101_io_in = _T_959 & io_rPort_8_en_0; // @[package.scala 94:16:@15113.4]
  assign RetimeWrapper_102_clock = clock; // @[:@15119.4]
  assign RetimeWrapper_102_reset = reset; // @[:@15120.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15122.4]
  assign RetimeWrapper_102_io_in = _T_1051 & io_rPort_8_en_0; // @[package.scala 94:16:@15121.4]
  assign RetimeWrapper_103_clock = clock; // @[:@15127.4]
  assign RetimeWrapper_103_reset = reset; // @[:@15128.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15130.4]
  assign RetimeWrapper_103_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@15129.4]
  assign RetimeWrapper_104_clock = clock; // @[:@15135.4]
  assign RetimeWrapper_104_reset = reset; // @[:@15136.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15138.4]
  assign RetimeWrapper_104_io_in = _T_1235 & io_rPort_8_en_0; // @[package.scala 94:16:@15137.4]
  assign RetimeWrapper_105_clock = clock; // @[:@15143.4]
  assign RetimeWrapper_105_reset = reset; // @[:@15144.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15146.4]
  assign RetimeWrapper_105_io_in = _T_1327 & io_rPort_8_en_0; // @[package.scala 94:16:@15145.4]
  assign RetimeWrapper_106_clock = clock; // @[:@15151.4]
  assign RetimeWrapper_106_reset = reset; // @[:@15152.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15154.4]
  assign RetimeWrapper_106_io_in = _T_1419 & io_rPort_8_en_0; // @[package.scala 94:16:@15153.4]
  assign RetimeWrapper_107_clock = clock; // @[:@15159.4]
  assign RetimeWrapper_107_reset = reset; // @[:@15160.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15162.4]
  assign RetimeWrapper_107_io_in = _T_1511 & io_rPort_8_en_0; // @[package.scala 94:16:@15161.4]
endmodule
module StickySelects_13( // @[:@16462.2]
  input   clock, // @[:@16463.4]
  input   reset, // @[:@16464.4]
  input   io_ins_0, // @[:@16465.4]
  input   io_ins_1, // @[:@16465.4]
  input   io_ins_2, // @[:@16465.4]
  input   io_ins_3, // @[:@16465.4]
  output  io_outs_0, // @[:@16465.4]
  output  io_outs_1, // @[:@16465.4]
  output  io_outs_2, // @[:@16465.4]
  output  io_outs_3 // @[:@16465.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@16467.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@16468.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@16469.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@16470.4]
  reg [31:0] _RAND_3;
  wire  _T_29; // @[StickySelects.scala 47:46:@16471.4]
  wire  _T_30; // @[StickySelects.scala 47:46:@16472.4]
  wire  _T_31; // @[StickySelects.scala 49:53:@16473.4]
  wire  _T_32; // @[StickySelects.scala 49:21:@16474.4]
  wire  _T_33; // @[StickySelects.scala 47:46:@16476.4]
  wire  _T_34; // @[StickySelects.scala 47:46:@16477.4]
  wire  _T_35; // @[StickySelects.scala 49:53:@16478.4]
  wire  _T_36; // @[StickySelects.scala 49:21:@16479.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@16481.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@16482.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@16483.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@16484.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@16487.4]
  wire  _T_43; // @[StickySelects.scala 49:53:@16488.4]
  wire  _T_44; // @[StickySelects.scala 49:21:@16489.4]
  assign _T_29 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@16471.4]
  assign _T_30 = _T_29 | io_ins_3; // @[StickySelects.scala 47:46:@16472.4]
  assign _T_31 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@16473.4]
  assign _T_32 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 49:21:@16474.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@16476.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 47:46:@16477.4]
  assign _T_35 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@16478.4]
  assign _T_36 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 49:21:@16479.4]
  assign _T_37 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@16481.4]
  assign _T_38 = _T_37 | io_ins_3; // @[StickySelects.scala 47:46:@16482.4]
  assign _T_39 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@16483.4]
  assign _T_40 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 49:21:@16484.4]
  assign _T_42 = _T_37 | io_ins_2; // @[StickySelects.scala 47:46:@16487.4]
  assign _T_43 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@16488.4]
  assign _T_44 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 49:21:@16489.4]
  assign io_outs_0 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 53:57:@16491.4]
  assign io_outs_1 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 53:57:@16492.4]
  assign io_outs_2 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 53:57:@16493.4]
  assign io_outs_3 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 53:57:@16494.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_30) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_31;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_35;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_39;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_42) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_43;
      end
    end
  end
endmodule
module x234_lb2_0( // @[:@18406.2]
  input         clock, // @[:@18407.4]
  input         reset, // @[:@18408.4]
  input  [1:0]  io_rPort_3_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_3_ofs_0, // @[:@18409.4]
  input         io_rPort_3_en_0, // @[:@18409.4]
  input         io_rPort_3_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_3_output_0, // @[:@18409.4]
  input  [1:0]  io_rPort_2_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_2_ofs_0, // @[:@18409.4]
  input         io_rPort_2_en_0, // @[:@18409.4]
  input         io_rPort_2_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_2_output_0, // @[:@18409.4]
  input  [1:0]  io_rPort_1_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_1_ofs_0, // @[:@18409.4]
  input         io_rPort_1_en_0, // @[:@18409.4]
  input         io_rPort_1_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_1_output_0, // @[:@18409.4]
  input  [1:0]  io_rPort_0_banks_1, // @[:@18409.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@18409.4]
  input  [9:0]  io_rPort_0_ofs_0, // @[:@18409.4]
  input         io_rPort_0_en_0, // @[:@18409.4]
  input         io_rPort_0_backpressure, // @[:@18409.4]
  output [31:0] io_rPort_0_output_0, // @[:@18409.4]
  input  [1:0]  io_wPort_0_banks_1, // @[:@18409.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@18409.4]
  input  [9:0]  io_wPort_0_ofs_0, // @[:@18409.4]
  input  [31:0] io_wPort_0_data_0, // @[:@18409.4]
  input         io_wPort_0_en_0 // @[:@18409.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [9:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [9:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@18444.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@18444.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [9:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [9:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@18460.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@18460.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [9:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [9:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@18476.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@18476.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [9:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [9:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@18492.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@18492.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [9:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [9:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@18508.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@18508.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [9:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [9:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@18524.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@18524.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [9:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [9:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@18540.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@18540.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [9:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [9:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@18556.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@18556.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [9:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [9:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@18572.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@18572.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [9:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [9:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@18588.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@18588.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [9:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [9:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@18604.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@18604.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [9:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [9:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@18620.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@18620.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@18796.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@18840.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@18884.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@18928.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@18972.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@19016.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@19060.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@19104.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@19148.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@19192.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@19236.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@19280.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@19345.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@19353.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@19361.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@19369.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@19377.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@19385.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@19393.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@19401.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@19409.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@19417.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@19425.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@19433.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@19489.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@19497.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@19505.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@19513.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@19521.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@19529.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@19537.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@19545.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@19553.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@19561.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@19569.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@19577.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@19633.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@19641.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@19649.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@19657.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@19665.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@19673.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@19681.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@19689.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@19697.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@19705.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@19713.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@19721.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@19777.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@19785.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@19793.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@19801.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@19809.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@19817.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@19825.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@19833.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@19841.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@19849.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@19857.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@19865.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@19865.4]
  wire  _T_166; // @[MemPrimitives.scala 82:210:@18636.4]
  wire  _T_168; // @[MemPrimitives.scala 82:210:@18637.4]
  wire  _T_169; // @[MemPrimitives.scala 82:228:@18638.4]
  wire  _T_170; // @[MemPrimitives.scala 83:102:@18639.4]
  wire [42:0] _T_172; // @[Cat.scala 30:58:@18641.4]
  wire  _T_179; // @[MemPrimitives.scala 82:210:@18649.4]
  wire  _T_180; // @[MemPrimitives.scala 82:228:@18650.4]
  wire  _T_181; // @[MemPrimitives.scala 83:102:@18651.4]
  wire [42:0] _T_183; // @[Cat.scala 30:58:@18653.4]
  wire  _T_190; // @[MemPrimitives.scala 82:210:@18661.4]
  wire  _T_191; // @[MemPrimitives.scala 82:228:@18662.4]
  wire  _T_192; // @[MemPrimitives.scala 83:102:@18663.4]
  wire [42:0] _T_194; // @[Cat.scala 30:58:@18665.4]
  wire  _T_199; // @[MemPrimitives.scala 82:210:@18672.4]
  wire  _T_202; // @[MemPrimitives.scala 82:228:@18674.4]
  wire  _T_203; // @[MemPrimitives.scala 83:102:@18675.4]
  wire [42:0] _T_205; // @[Cat.scala 30:58:@18677.4]
  wire  _T_213; // @[MemPrimitives.scala 82:228:@18686.4]
  wire  _T_214; // @[MemPrimitives.scala 83:102:@18687.4]
  wire [42:0] _T_216; // @[Cat.scala 30:58:@18689.4]
  wire  _T_224; // @[MemPrimitives.scala 82:228:@18698.4]
  wire  _T_225; // @[MemPrimitives.scala 83:102:@18699.4]
  wire [42:0] _T_227; // @[Cat.scala 30:58:@18701.4]
  wire  _T_232; // @[MemPrimitives.scala 82:210:@18708.4]
  wire  _T_235; // @[MemPrimitives.scala 82:228:@18710.4]
  wire  _T_236; // @[MemPrimitives.scala 83:102:@18711.4]
  wire [42:0] _T_238; // @[Cat.scala 30:58:@18713.4]
  wire  _T_246; // @[MemPrimitives.scala 82:228:@18722.4]
  wire  _T_247; // @[MemPrimitives.scala 83:102:@18723.4]
  wire [42:0] _T_249; // @[Cat.scala 30:58:@18725.4]
  wire  _T_257; // @[MemPrimitives.scala 82:228:@18734.4]
  wire  _T_258; // @[MemPrimitives.scala 83:102:@18735.4]
  wire [42:0] _T_260; // @[Cat.scala 30:58:@18737.4]
  wire  _T_265; // @[MemPrimitives.scala 82:210:@18744.4]
  wire  _T_268; // @[MemPrimitives.scala 82:228:@18746.4]
  wire  _T_269; // @[MemPrimitives.scala 83:102:@18747.4]
  wire [42:0] _T_271; // @[Cat.scala 30:58:@18749.4]
  wire  _T_279; // @[MemPrimitives.scala 82:228:@18758.4]
  wire  _T_280; // @[MemPrimitives.scala 83:102:@18759.4]
  wire [42:0] _T_282; // @[Cat.scala 30:58:@18761.4]
  wire  _T_290; // @[MemPrimitives.scala 82:228:@18770.4]
  wire  _T_291; // @[MemPrimitives.scala 83:102:@18771.4]
  wire [42:0] _T_293; // @[Cat.scala 30:58:@18773.4]
  wire  _T_298; // @[MemPrimitives.scala 110:210:@18780.4]
  wire  _T_300; // @[MemPrimitives.scala 110:210:@18781.4]
  wire  _T_301; // @[MemPrimitives.scala 110:228:@18782.4]
  wire  _T_304; // @[MemPrimitives.scala 110:210:@18784.4]
  wire  _T_306; // @[MemPrimitives.scala 110:210:@18785.4]
  wire  _T_307; // @[MemPrimitives.scala 110:228:@18786.4]
  wire  _T_310; // @[MemPrimitives.scala 110:210:@18788.4]
  wire  _T_312; // @[MemPrimitives.scala 110:210:@18789.4]
  wire  _T_313; // @[MemPrimitives.scala 110:228:@18790.4]
  wire  _T_316; // @[MemPrimitives.scala 110:210:@18792.4]
  wire  _T_318; // @[MemPrimitives.scala 110:210:@18793.4]
  wire  _T_319; // @[MemPrimitives.scala 110:228:@18794.4]
  wire  _T_321; // @[MemPrimitives.scala 126:35:@18803.4]
  wire  _T_322; // @[MemPrimitives.scala 126:35:@18804.4]
  wire  _T_323; // @[MemPrimitives.scala 126:35:@18805.4]
  wire  _T_324; // @[MemPrimitives.scala 126:35:@18806.4]
  wire [11:0] _T_326; // @[Cat.scala 30:58:@18808.4]
  wire [11:0] _T_328; // @[Cat.scala 30:58:@18810.4]
  wire [11:0] _T_330; // @[Cat.scala 30:58:@18812.4]
  wire [11:0] _T_332; // @[Cat.scala 30:58:@18814.4]
  wire [11:0] _T_333; // @[Mux.scala 31:69:@18815.4]
  wire [11:0] _T_334; // @[Mux.scala 31:69:@18816.4]
  wire [11:0] _T_335; // @[Mux.scala 31:69:@18817.4]
  wire  _T_342; // @[MemPrimitives.scala 110:210:@18825.4]
  wire  _T_343; // @[MemPrimitives.scala 110:228:@18826.4]
  wire  _T_348; // @[MemPrimitives.scala 110:210:@18829.4]
  wire  _T_349; // @[MemPrimitives.scala 110:228:@18830.4]
  wire  _T_354; // @[MemPrimitives.scala 110:210:@18833.4]
  wire  _T_355; // @[MemPrimitives.scala 110:228:@18834.4]
  wire  _T_360; // @[MemPrimitives.scala 110:210:@18837.4]
  wire  _T_361; // @[MemPrimitives.scala 110:228:@18838.4]
  wire  _T_363; // @[MemPrimitives.scala 126:35:@18847.4]
  wire  _T_364; // @[MemPrimitives.scala 126:35:@18848.4]
  wire  _T_365; // @[MemPrimitives.scala 126:35:@18849.4]
  wire  _T_366; // @[MemPrimitives.scala 126:35:@18850.4]
  wire [11:0] _T_368; // @[Cat.scala 30:58:@18852.4]
  wire [11:0] _T_370; // @[Cat.scala 30:58:@18854.4]
  wire [11:0] _T_372; // @[Cat.scala 30:58:@18856.4]
  wire [11:0] _T_374; // @[Cat.scala 30:58:@18858.4]
  wire [11:0] _T_375; // @[Mux.scala 31:69:@18859.4]
  wire [11:0] _T_376; // @[Mux.scala 31:69:@18860.4]
  wire [11:0] _T_377; // @[Mux.scala 31:69:@18861.4]
  wire  _T_384; // @[MemPrimitives.scala 110:210:@18869.4]
  wire  _T_385; // @[MemPrimitives.scala 110:228:@18870.4]
  wire  _T_390; // @[MemPrimitives.scala 110:210:@18873.4]
  wire  _T_391; // @[MemPrimitives.scala 110:228:@18874.4]
  wire  _T_396; // @[MemPrimitives.scala 110:210:@18877.4]
  wire  _T_397; // @[MemPrimitives.scala 110:228:@18878.4]
  wire  _T_402; // @[MemPrimitives.scala 110:210:@18881.4]
  wire  _T_403; // @[MemPrimitives.scala 110:228:@18882.4]
  wire  _T_405; // @[MemPrimitives.scala 126:35:@18891.4]
  wire  _T_406; // @[MemPrimitives.scala 126:35:@18892.4]
  wire  _T_407; // @[MemPrimitives.scala 126:35:@18893.4]
  wire  _T_408; // @[MemPrimitives.scala 126:35:@18894.4]
  wire [11:0] _T_410; // @[Cat.scala 30:58:@18896.4]
  wire [11:0] _T_412; // @[Cat.scala 30:58:@18898.4]
  wire [11:0] _T_414; // @[Cat.scala 30:58:@18900.4]
  wire [11:0] _T_416; // @[Cat.scala 30:58:@18902.4]
  wire [11:0] _T_417; // @[Mux.scala 31:69:@18903.4]
  wire [11:0] _T_418; // @[Mux.scala 31:69:@18904.4]
  wire [11:0] _T_419; // @[Mux.scala 31:69:@18905.4]
  wire  _T_424; // @[MemPrimitives.scala 110:210:@18912.4]
  wire  _T_427; // @[MemPrimitives.scala 110:228:@18914.4]
  wire  _T_430; // @[MemPrimitives.scala 110:210:@18916.4]
  wire  _T_433; // @[MemPrimitives.scala 110:228:@18918.4]
  wire  _T_436; // @[MemPrimitives.scala 110:210:@18920.4]
  wire  _T_439; // @[MemPrimitives.scala 110:228:@18922.4]
  wire  _T_442; // @[MemPrimitives.scala 110:210:@18924.4]
  wire  _T_445; // @[MemPrimitives.scala 110:228:@18926.4]
  wire  _T_447; // @[MemPrimitives.scala 126:35:@18935.4]
  wire  _T_448; // @[MemPrimitives.scala 126:35:@18936.4]
  wire  _T_449; // @[MemPrimitives.scala 126:35:@18937.4]
  wire  _T_450; // @[MemPrimitives.scala 126:35:@18938.4]
  wire [11:0] _T_452; // @[Cat.scala 30:58:@18940.4]
  wire [11:0] _T_454; // @[Cat.scala 30:58:@18942.4]
  wire [11:0] _T_456; // @[Cat.scala 30:58:@18944.4]
  wire [11:0] _T_458; // @[Cat.scala 30:58:@18946.4]
  wire [11:0] _T_459; // @[Mux.scala 31:69:@18947.4]
  wire [11:0] _T_460; // @[Mux.scala 31:69:@18948.4]
  wire [11:0] _T_461; // @[Mux.scala 31:69:@18949.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@18958.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@18962.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@18966.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@18970.4]
  wire  _T_489; // @[MemPrimitives.scala 126:35:@18979.4]
  wire  _T_490; // @[MemPrimitives.scala 126:35:@18980.4]
  wire  _T_491; // @[MemPrimitives.scala 126:35:@18981.4]
  wire  _T_492; // @[MemPrimitives.scala 126:35:@18982.4]
  wire [11:0] _T_494; // @[Cat.scala 30:58:@18984.4]
  wire [11:0] _T_496; // @[Cat.scala 30:58:@18986.4]
  wire [11:0] _T_498; // @[Cat.scala 30:58:@18988.4]
  wire [11:0] _T_500; // @[Cat.scala 30:58:@18990.4]
  wire [11:0] _T_501; // @[Mux.scala 31:69:@18991.4]
  wire [11:0] _T_502; // @[Mux.scala 31:69:@18992.4]
  wire [11:0] _T_503; // @[Mux.scala 31:69:@18993.4]
  wire  _T_511; // @[MemPrimitives.scala 110:228:@19002.4]
  wire  _T_517; // @[MemPrimitives.scala 110:228:@19006.4]
  wire  _T_523; // @[MemPrimitives.scala 110:228:@19010.4]
  wire  _T_529; // @[MemPrimitives.scala 110:228:@19014.4]
  wire  _T_531; // @[MemPrimitives.scala 126:35:@19023.4]
  wire  _T_532; // @[MemPrimitives.scala 126:35:@19024.4]
  wire  _T_533; // @[MemPrimitives.scala 126:35:@19025.4]
  wire  _T_534; // @[MemPrimitives.scala 126:35:@19026.4]
  wire [11:0] _T_536; // @[Cat.scala 30:58:@19028.4]
  wire [11:0] _T_538; // @[Cat.scala 30:58:@19030.4]
  wire [11:0] _T_540; // @[Cat.scala 30:58:@19032.4]
  wire [11:0] _T_542; // @[Cat.scala 30:58:@19034.4]
  wire [11:0] _T_543; // @[Mux.scala 31:69:@19035.4]
  wire [11:0] _T_544; // @[Mux.scala 31:69:@19036.4]
  wire [11:0] _T_545; // @[Mux.scala 31:69:@19037.4]
  wire  _T_550; // @[MemPrimitives.scala 110:210:@19044.4]
  wire  _T_553; // @[MemPrimitives.scala 110:228:@19046.4]
  wire  _T_556; // @[MemPrimitives.scala 110:210:@19048.4]
  wire  _T_559; // @[MemPrimitives.scala 110:228:@19050.4]
  wire  _T_562; // @[MemPrimitives.scala 110:210:@19052.4]
  wire  _T_565; // @[MemPrimitives.scala 110:228:@19054.4]
  wire  _T_568; // @[MemPrimitives.scala 110:210:@19056.4]
  wire  _T_571; // @[MemPrimitives.scala 110:228:@19058.4]
  wire  _T_573; // @[MemPrimitives.scala 126:35:@19067.4]
  wire  _T_574; // @[MemPrimitives.scala 126:35:@19068.4]
  wire  _T_575; // @[MemPrimitives.scala 126:35:@19069.4]
  wire  _T_576; // @[MemPrimitives.scala 126:35:@19070.4]
  wire [11:0] _T_578; // @[Cat.scala 30:58:@19072.4]
  wire [11:0] _T_580; // @[Cat.scala 30:58:@19074.4]
  wire [11:0] _T_582; // @[Cat.scala 30:58:@19076.4]
  wire [11:0] _T_584; // @[Cat.scala 30:58:@19078.4]
  wire [11:0] _T_585; // @[Mux.scala 31:69:@19079.4]
  wire [11:0] _T_586; // @[Mux.scala 31:69:@19080.4]
  wire [11:0] _T_587; // @[Mux.scala 31:69:@19081.4]
  wire  _T_595; // @[MemPrimitives.scala 110:228:@19090.4]
  wire  _T_601; // @[MemPrimitives.scala 110:228:@19094.4]
  wire  _T_607; // @[MemPrimitives.scala 110:228:@19098.4]
  wire  _T_613; // @[MemPrimitives.scala 110:228:@19102.4]
  wire  _T_615; // @[MemPrimitives.scala 126:35:@19111.4]
  wire  _T_616; // @[MemPrimitives.scala 126:35:@19112.4]
  wire  _T_617; // @[MemPrimitives.scala 126:35:@19113.4]
  wire  _T_618; // @[MemPrimitives.scala 126:35:@19114.4]
  wire [11:0] _T_620; // @[Cat.scala 30:58:@19116.4]
  wire [11:0] _T_622; // @[Cat.scala 30:58:@19118.4]
  wire [11:0] _T_624; // @[Cat.scala 30:58:@19120.4]
  wire [11:0] _T_626; // @[Cat.scala 30:58:@19122.4]
  wire [11:0] _T_627; // @[Mux.scala 31:69:@19123.4]
  wire [11:0] _T_628; // @[Mux.scala 31:69:@19124.4]
  wire [11:0] _T_629; // @[Mux.scala 31:69:@19125.4]
  wire  _T_637; // @[MemPrimitives.scala 110:228:@19134.4]
  wire  _T_643; // @[MemPrimitives.scala 110:228:@19138.4]
  wire  _T_649; // @[MemPrimitives.scala 110:228:@19142.4]
  wire  _T_655; // @[MemPrimitives.scala 110:228:@19146.4]
  wire  _T_657; // @[MemPrimitives.scala 126:35:@19155.4]
  wire  _T_658; // @[MemPrimitives.scala 126:35:@19156.4]
  wire  _T_659; // @[MemPrimitives.scala 126:35:@19157.4]
  wire  _T_660; // @[MemPrimitives.scala 126:35:@19158.4]
  wire [11:0] _T_662; // @[Cat.scala 30:58:@19160.4]
  wire [11:0] _T_664; // @[Cat.scala 30:58:@19162.4]
  wire [11:0] _T_666; // @[Cat.scala 30:58:@19164.4]
  wire [11:0] _T_668; // @[Cat.scala 30:58:@19166.4]
  wire [11:0] _T_669; // @[Mux.scala 31:69:@19167.4]
  wire [11:0] _T_670; // @[Mux.scala 31:69:@19168.4]
  wire [11:0] _T_671; // @[Mux.scala 31:69:@19169.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@19176.4]
  wire  _T_679; // @[MemPrimitives.scala 110:228:@19178.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@19180.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@19182.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@19184.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@19186.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@19188.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@19190.4]
  wire  _T_699; // @[MemPrimitives.scala 126:35:@19199.4]
  wire  _T_700; // @[MemPrimitives.scala 126:35:@19200.4]
  wire  _T_701; // @[MemPrimitives.scala 126:35:@19201.4]
  wire  _T_702; // @[MemPrimitives.scala 126:35:@19202.4]
  wire [11:0] _T_704; // @[Cat.scala 30:58:@19204.4]
  wire [11:0] _T_706; // @[Cat.scala 30:58:@19206.4]
  wire [11:0] _T_708; // @[Cat.scala 30:58:@19208.4]
  wire [11:0] _T_710; // @[Cat.scala 30:58:@19210.4]
  wire [11:0] _T_711; // @[Mux.scala 31:69:@19211.4]
  wire [11:0] _T_712; // @[Mux.scala 31:69:@19212.4]
  wire [11:0] _T_713; // @[Mux.scala 31:69:@19213.4]
  wire  _T_721; // @[MemPrimitives.scala 110:228:@19222.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@19226.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@19230.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@19234.4]
  wire  _T_741; // @[MemPrimitives.scala 126:35:@19243.4]
  wire  _T_742; // @[MemPrimitives.scala 126:35:@19244.4]
  wire  _T_743; // @[MemPrimitives.scala 126:35:@19245.4]
  wire  _T_744; // @[MemPrimitives.scala 126:35:@19246.4]
  wire [11:0] _T_746; // @[Cat.scala 30:58:@19248.4]
  wire [11:0] _T_748; // @[Cat.scala 30:58:@19250.4]
  wire [11:0] _T_750; // @[Cat.scala 30:58:@19252.4]
  wire [11:0] _T_752; // @[Cat.scala 30:58:@19254.4]
  wire [11:0] _T_753; // @[Mux.scala 31:69:@19255.4]
  wire [11:0] _T_754; // @[Mux.scala 31:69:@19256.4]
  wire [11:0] _T_755; // @[Mux.scala 31:69:@19257.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@19266.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@19270.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@19274.4]
  wire  _T_781; // @[MemPrimitives.scala 110:228:@19278.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@19287.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@19288.4]
  wire  _T_785; // @[MemPrimitives.scala 126:35:@19289.4]
  wire  _T_786; // @[MemPrimitives.scala 126:35:@19290.4]
  wire [11:0] _T_788; // @[Cat.scala 30:58:@19292.4]
  wire [11:0] _T_790; // @[Cat.scala 30:58:@19294.4]
  wire [11:0] _T_792; // @[Cat.scala 30:58:@19296.4]
  wire [11:0] _T_794; // @[Cat.scala 30:58:@19298.4]
  wire [11:0] _T_795; // @[Mux.scala 31:69:@19299.4]
  wire [11:0] _T_796; // @[Mux.scala 31:69:@19300.4]
  wire [11:0] _T_797; // @[Mux.scala 31:69:@19301.4]
  wire  _T_893; // @[package.scala 96:25:@19430.4 package.scala 96:25:@19431.4]
  wire [31:0] _T_897; // @[Mux.scala 31:69:@19440.4]
  wire  _T_890; // @[package.scala 96:25:@19422.4 package.scala 96:25:@19423.4]
  wire [31:0] _T_898; // @[Mux.scala 31:69:@19441.4]
  wire  _T_887; // @[package.scala 96:25:@19414.4 package.scala 96:25:@19415.4]
  wire [31:0] _T_899; // @[Mux.scala 31:69:@19442.4]
  wire  _T_884; // @[package.scala 96:25:@19406.4 package.scala 96:25:@19407.4]
  wire [31:0] _T_900; // @[Mux.scala 31:69:@19443.4]
  wire  _T_881; // @[package.scala 96:25:@19398.4 package.scala 96:25:@19399.4]
  wire [31:0] _T_901; // @[Mux.scala 31:69:@19444.4]
  wire  _T_878; // @[package.scala 96:25:@19390.4 package.scala 96:25:@19391.4]
  wire [31:0] _T_902; // @[Mux.scala 31:69:@19445.4]
  wire  _T_875; // @[package.scala 96:25:@19382.4 package.scala 96:25:@19383.4]
  wire [31:0] _T_903; // @[Mux.scala 31:69:@19446.4]
  wire  _T_872; // @[package.scala 96:25:@19374.4 package.scala 96:25:@19375.4]
  wire [31:0] _T_904; // @[Mux.scala 31:69:@19447.4]
  wire  _T_869; // @[package.scala 96:25:@19366.4 package.scala 96:25:@19367.4]
  wire [31:0] _T_905; // @[Mux.scala 31:69:@19448.4]
  wire  _T_866; // @[package.scala 96:25:@19358.4 package.scala 96:25:@19359.4]
  wire [31:0] _T_906; // @[Mux.scala 31:69:@19449.4]
  wire  _T_863; // @[package.scala 96:25:@19350.4 package.scala 96:25:@19351.4]
  wire  _T_1000; // @[package.scala 96:25:@19574.4 package.scala 96:25:@19575.4]
  wire [31:0] _T_1004; // @[Mux.scala 31:69:@19584.4]
  wire  _T_997; // @[package.scala 96:25:@19566.4 package.scala 96:25:@19567.4]
  wire [31:0] _T_1005; // @[Mux.scala 31:69:@19585.4]
  wire  _T_994; // @[package.scala 96:25:@19558.4 package.scala 96:25:@19559.4]
  wire [31:0] _T_1006; // @[Mux.scala 31:69:@19586.4]
  wire  _T_991; // @[package.scala 96:25:@19550.4 package.scala 96:25:@19551.4]
  wire [31:0] _T_1007; // @[Mux.scala 31:69:@19587.4]
  wire  _T_988; // @[package.scala 96:25:@19542.4 package.scala 96:25:@19543.4]
  wire [31:0] _T_1008; // @[Mux.scala 31:69:@19588.4]
  wire  _T_985; // @[package.scala 96:25:@19534.4 package.scala 96:25:@19535.4]
  wire [31:0] _T_1009; // @[Mux.scala 31:69:@19589.4]
  wire  _T_982; // @[package.scala 96:25:@19526.4 package.scala 96:25:@19527.4]
  wire [31:0] _T_1010; // @[Mux.scala 31:69:@19590.4]
  wire  _T_979; // @[package.scala 96:25:@19518.4 package.scala 96:25:@19519.4]
  wire [31:0] _T_1011; // @[Mux.scala 31:69:@19591.4]
  wire  _T_976; // @[package.scala 96:25:@19510.4 package.scala 96:25:@19511.4]
  wire [31:0] _T_1012; // @[Mux.scala 31:69:@19592.4]
  wire  _T_973; // @[package.scala 96:25:@19502.4 package.scala 96:25:@19503.4]
  wire [31:0] _T_1013; // @[Mux.scala 31:69:@19593.4]
  wire  _T_970; // @[package.scala 96:25:@19494.4 package.scala 96:25:@19495.4]
  wire  _T_1107; // @[package.scala 96:25:@19718.4 package.scala 96:25:@19719.4]
  wire [31:0] _T_1111; // @[Mux.scala 31:69:@19728.4]
  wire  _T_1104; // @[package.scala 96:25:@19710.4 package.scala 96:25:@19711.4]
  wire [31:0] _T_1112; // @[Mux.scala 31:69:@19729.4]
  wire  _T_1101; // @[package.scala 96:25:@19702.4 package.scala 96:25:@19703.4]
  wire [31:0] _T_1113; // @[Mux.scala 31:69:@19730.4]
  wire  _T_1098; // @[package.scala 96:25:@19694.4 package.scala 96:25:@19695.4]
  wire [31:0] _T_1114; // @[Mux.scala 31:69:@19731.4]
  wire  _T_1095; // @[package.scala 96:25:@19686.4 package.scala 96:25:@19687.4]
  wire [31:0] _T_1115; // @[Mux.scala 31:69:@19732.4]
  wire  _T_1092; // @[package.scala 96:25:@19678.4 package.scala 96:25:@19679.4]
  wire [31:0] _T_1116; // @[Mux.scala 31:69:@19733.4]
  wire  _T_1089; // @[package.scala 96:25:@19670.4 package.scala 96:25:@19671.4]
  wire [31:0] _T_1117; // @[Mux.scala 31:69:@19734.4]
  wire  _T_1086; // @[package.scala 96:25:@19662.4 package.scala 96:25:@19663.4]
  wire [31:0] _T_1118; // @[Mux.scala 31:69:@19735.4]
  wire  _T_1083; // @[package.scala 96:25:@19654.4 package.scala 96:25:@19655.4]
  wire [31:0] _T_1119; // @[Mux.scala 31:69:@19736.4]
  wire  _T_1080; // @[package.scala 96:25:@19646.4 package.scala 96:25:@19647.4]
  wire [31:0] _T_1120; // @[Mux.scala 31:69:@19737.4]
  wire  _T_1077; // @[package.scala 96:25:@19638.4 package.scala 96:25:@19639.4]
  wire  _T_1214; // @[package.scala 96:25:@19862.4 package.scala 96:25:@19863.4]
  wire [31:0] _T_1218; // @[Mux.scala 31:69:@19872.4]
  wire  _T_1211; // @[package.scala 96:25:@19854.4 package.scala 96:25:@19855.4]
  wire [31:0] _T_1219; // @[Mux.scala 31:69:@19873.4]
  wire  _T_1208; // @[package.scala 96:25:@19846.4 package.scala 96:25:@19847.4]
  wire [31:0] _T_1220; // @[Mux.scala 31:69:@19874.4]
  wire  _T_1205; // @[package.scala 96:25:@19838.4 package.scala 96:25:@19839.4]
  wire [31:0] _T_1221; // @[Mux.scala 31:69:@19875.4]
  wire  _T_1202; // @[package.scala 96:25:@19830.4 package.scala 96:25:@19831.4]
  wire [31:0] _T_1222; // @[Mux.scala 31:69:@19876.4]
  wire  _T_1199; // @[package.scala 96:25:@19822.4 package.scala 96:25:@19823.4]
  wire [31:0] _T_1223; // @[Mux.scala 31:69:@19877.4]
  wire  _T_1196; // @[package.scala 96:25:@19814.4 package.scala 96:25:@19815.4]
  wire [31:0] _T_1224; // @[Mux.scala 31:69:@19878.4]
  wire  _T_1193; // @[package.scala 96:25:@19806.4 package.scala 96:25:@19807.4]
  wire [31:0] _T_1225; // @[Mux.scala 31:69:@19879.4]
  wire  _T_1190; // @[package.scala 96:25:@19798.4 package.scala 96:25:@19799.4]
  wire [31:0] _T_1226; // @[Mux.scala 31:69:@19880.4]
  wire  _T_1187; // @[package.scala 96:25:@19790.4 package.scala 96:25:@19791.4]
  wire [31:0] _T_1227; // @[Mux.scala 31:69:@19881.4]
  wire  _T_1184; // @[package.scala 96:25:@19782.4 package.scala 96:25:@19783.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@18444.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@18460.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@18476.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@18492.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@18508.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@18524.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@18540.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@18556.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@18572.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@18588.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@18604.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@18620.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects_13 StickySelects ( // @[MemPrimitives.scala 124:33:@18796.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3)
  );
  StickySelects_13 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@18840.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_13 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@18884.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3)
  );
  StickySelects_13 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@18928.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3)
  );
  StickySelects_13 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@18972.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3)
  );
  StickySelects_13 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@19016.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_13 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@19060.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3)
  );
  StickySelects_13 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@19104.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3)
  );
  StickySelects_13 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@19148.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3)
  );
  StickySelects_13 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@19192.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_13 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@19236.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3)
  );
  StickySelects_13 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@19280.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@19345.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@19353.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@19361.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@19369.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@19377.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@19385.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@19393.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@19401.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@19409.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@19417.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@19425.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@19433.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@19489.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@19497.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@19505.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@19513.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@19521.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@19529.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@19537.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@19545.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@19553.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@19561.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@19569.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@19577.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@19633.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@19641.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@19649.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@19657.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@19665.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@19673.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@19681.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@19689.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@19697.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@19705.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@19713.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@19721.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@19777.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@19785.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@19793.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@19801.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@19809.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@19817.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@19825.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@19833.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@19841.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@19849.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@19857.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@19865.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  assign _T_166 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@18636.4]
  assign _T_168 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@18637.4]
  assign _T_169 = _T_166 & _T_168; // @[MemPrimitives.scala 82:228:@18638.4]
  assign _T_170 = io_wPort_0_en_0 & _T_169; // @[MemPrimitives.scala 83:102:@18639.4]
  assign _T_172 = {_T_170,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18641.4]
  assign _T_179 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@18649.4]
  assign _T_180 = _T_166 & _T_179; // @[MemPrimitives.scala 82:228:@18650.4]
  assign _T_181 = io_wPort_0_en_0 & _T_180; // @[MemPrimitives.scala 83:102:@18651.4]
  assign _T_183 = {_T_181,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18653.4]
  assign _T_190 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@18661.4]
  assign _T_191 = _T_166 & _T_190; // @[MemPrimitives.scala 82:228:@18662.4]
  assign _T_192 = io_wPort_0_en_0 & _T_191; // @[MemPrimitives.scala 83:102:@18663.4]
  assign _T_194 = {_T_192,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18665.4]
  assign _T_199 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@18672.4]
  assign _T_202 = _T_199 & _T_168; // @[MemPrimitives.scala 82:228:@18674.4]
  assign _T_203 = io_wPort_0_en_0 & _T_202; // @[MemPrimitives.scala 83:102:@18675.4]
  assign _T_205 = {_T_203,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18677.4]
  assign _T_213 = _T_199 & _T_179; // @[MemPrimitives.scala 82:228:@18686.4]
  assign _T_214 = io_wPort_0_en_0 & _T_213; // @[MemPrimitives.scala 83:102:@18687.4]
  assign _T_216 = {_T_214,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18689.4]
  assign _T_224 = _T_199 & _T_190; // @[MemPrimitives.scala 82:228:@18698.4]
  assign _T_225 = io_wPort_0_en_0 & _T_224; // @[MemPrimitives.scala 83:102:@18699.4]
  assign _T_227 = {_T_225,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18701.4]
  assign _T_232 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@18708.4]
  assign _T_235 = _T_232 & _T_168; // @[MemPrimitives.scala 82:228:@18710.4]
  assign _T_236 = io_wPort_0_en_0 & _T_235; // @[MemPrimitives.scala 83:102:@18711.4]
  assign _T_238 = {_T_236,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18713.4]
  assign _T_246 = _T_232 & _T_179; // @[MemPrimitives.scala 82:228:@18722.4]
  assign _T_247 = io_wPort_0_en_0 & _T_246; // @[MemPrimitives.scala 83:102:@18723.4]
  assign _T_249 = {_T_247,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18725.4]
  assign _T_257 = _T_232 & _T_190; // @[MemPrimitives.scala 82:228:@18734.4]
  assign _T_258 = io_wPort_0_en_0 & _T_257; // @[MemPrimitives.scala 83:102:@18735.4]
  assign _T_260 = {_T_258,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18737.4]
  assign _T_265 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@18744.4]
  assign _T_268 = _T_265 & _T_168; // @[MemPrimitives.scala 82:228:@18746.4]
  assign _T_269 = io_wPort_0_en_0 & _T_268; // @[MemPrimitives.scala 83:102:@18747.4]
  assign _T_271 = {_T_269,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18749.4]
  assign _T_279 = _T_265 & _T_179; // @[MemPrimitives.scala 82:228:@18758.4]
  assign _T_280 = io_wPort_0_en_0 & _T_279; // @[MemPrimitives.scala 83:102:@18759.4]
  assign _T_282 = {_T_280,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18761.4]
  assign _T_290 = _T_265 & _T_190; // @[MemPrimitives.scala 82:228:@18770.4]
  assign _T_291 = io_wPort_0_en_0 & _T_290; // @[MemPrimitives.scala 83:102:@18771.4]
  assign _T_293 = {_T_291,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18773.4]
  assign _T_298 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18780.4]
  assign _T_300 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18781.4]
  assign _T_301 = _T_298 & _T_300; // @[MemPrimitives.scala 110:228:@18782.4]
  assign _T_304 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18784.4]
  assign _T_306 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18785.4]
  assign _T_307 = _T_304 & _T_306; // @[MemPrimitives.scala 110:228:@18786.4]
  assign _T_310 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18788.4]
  assign _T_312 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18789.4]
  assign _T_313 = _T_310 & _T_312; // @[MemPrimitives.scala 110:228:@18790.4]
  assign _T_316 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@18792.4]
  assign _T_318 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@18793.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 110:228:@18794.4]
  assign _T_321 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@18803.4]
  assign _T_322 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@18804.4]
  assign _T_323 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@18805.4]
  assign _T_324 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@18806.4]
  assign _T_326 = {_T_321,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18808.4]
  assign _T_328 = {_T_322,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18810.4]
  assign _T_330 = {_T_323,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18812.4]
  assign _T_332 = {_T_324,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18814.4]
  assign _T_333 = _T_323 ? _T_330 : _T_332; // @[Mux.scala 31:69:@18815.4]
  assign _T_334 = _T_322 ? _T_328 : _T_333; // @[Mux.scala 31:69:@18816.4]
  assign _T_335 = _T_321 ? _T_326 : _T_334; // @[Mux.scala 31:69:@18817.4]
  assign _T_342 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18825.4]
  assign _T_343 = _T_298 & _T_342; // @[MemPrimitives.scala 110:228:@18826.4]
  assign _T_348 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18829.4]
  assign _T_349 = _T_304 & _T_348; // @[MemPrimitives.scala 110:228:@18830.4]
  assign _T_354 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18833.4]
  assign _T_355 = _T_310 & _T_354; // @[MemPrimitives.scala 110:228:@18834.4]
  assign _T_360 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@18837.4]
  assign _T_361 = _T_316 & _T_360; // @[MemPrimitives.scala 110:228:@18838.4]
  assign _T_363 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@18847.4]
  assign _T_364 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@18848.4]
  assign _T_365 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@18849.4]
  assign _T_366 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@18850.4]
  assign _T_368 = {_T_363,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18852.4]
  assign _T_370 = {_T_364,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18854.4]
  assign _T_372 = {_T_365,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18856.4]
  assign _T_374 = {_T_366,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18858.4]
  assign _T_375 = _T_365 ? _T_372 : _T_374; // @[Mux.scala 31:69:@18859.4]
  assign _T_376 = _T_364 ? _T_370 : _T_375; // @[Mux.scala 31:69:@18860.4]
  assign _T_377 = _T_363 ? _T_368 : _T_376; // @[Mux.scala 31:69:@18861.4]
  assign _T_384 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18869.4]
  assign _T_385 = _T_298 & _T_384; // @[MemPrimitives.scala 110:228:@18870.4]
  assign _T_390 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18873.4]
  assign _T_391 = _T_304 & _T_390; // @[MemPrimitives.scala 110:228:@18874.4]
  assign _T_396 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18877.4]
  assign _T_397 = _T_310 & _T_396; // @[MemPrimitives.scala 110:228:@18878.4]
  assign _T_402 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@18881.4]
  assign _T_403 = _T_316 & _T_402; // @[MemPrimitives.scala 110:228:@18882.4]
  assign _T_405 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@18891.4]
  assign _T_406 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@18892.4]
  assign _T_407 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@18893.4]
  assign _T_408 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@18894.4]
  assign _T_410 = {_T_405,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18896.4]
  assign _T_412 = {_T_406,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18898.4]
  assign _T_414 = {_T_407,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18900.4]
  assign _T_416 = {_T_408,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18902.4]
  assign _T_417 = _T_407 ? _T_414 : _T_416; // @[Mux.scala 31:69:@18903.4]
  assign _T_418 = _T_406 ? _T_412 : _T_417; // @[Mux.scala 31:69:@18904.4]
  assign _T_419 = _T_405 ? _T_410 : _T_418; // @[Mux.scala 31:69:@18905.4]
  assign _T_424 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18912.4]
  assign _T_427 = _T_424 & _T_300; // @[MemPrimitives.scala 110:228:@18914.4]
  assign _T_430 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18916.4]
  assign _T_433 = _T_430 & _T_306; // @[MemPrimitives.scala 110:228:@18918.4]
  assign _T_436 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18920.4]
  assign _T_439 = _T_436 & _T_312; // @[MemPrimitives.scala 110:228:@18922.4]
  assign _T_442 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@18924.4]
  assign _T_445 = _T_442 & _T_318; // @[MemPrimitives.scala 110:228:@18926.4]
  assign _T_447 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@18935.4]
  assign _T_448 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@18936.4]
  assign _T_449 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@18937.4]
  assign _T_450 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@18938.4]
  assign _T_452 = {_T_447,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18940.4]
  assign _T_454 = {_T_448,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18942.4]
  assign _T_456 = {_T_449,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18944.4]
  assign _T_458 = {_T_450,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18946.4]
  assign _T_459 = _T_449 ? _T_456 : _T_458; // @[Mux.scala 31:69:@18947.4]
  assign _T_460 = _T_448 ? _T_454 : _T_459; // @[Mux.scala 31:69:@18948.4]
  assign _T_461 = _T_447 ? _T_452 : _T_460; // @[Mux.scala 31:69:@18949.4]
  assign _T_469 = _T_424 & _T_342; // @[MemPrimitives.scala 110:228:@18958.4]
  assign _T_475 = _T_430 & _T_348; // @[MemPrimitives.scala 110:228:@18962.4]
  assign _T_481 = _T_436 & _T_354; // @[MemPrimitives.scala 110:228:@18966.4]
  assign _T_487 = _T_442 & _T_360; // @[MemPrimitives.scala 110:228:@18970.4]
  assign _T_489 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@18979.4]
  assign _T_490 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@18980.4]
  assign _T_491 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@18981.4]
  assign _T_492 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@18982.4]
  assign _T_494 = {_T_489,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@18984.4]
  assign _T_496 = {_T_490,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@18986.4]
  assign _T_498 = {_T_491,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@18988.4]
  assign _T_500 = {_T_492,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@18990.4]
  assign _T_501 = _T_491 ? _T_498 : _T_500; // @[Mux.scala 31:69:@18991.4]
  assign _T_502 = _T_490 ? _T_496 : _T_501; // @[Mux.scala 31:69:@18992.4]
  assign _T_503 = _T_489 ? _T_494 : _T_502; // @[Mux.scala 31:69:@18993.4]
  assign _T_511 = _T_424 & _T_384; // @[MemPrimitives.scala 110:228:@19002.4]
  assign _T_517 = _T_430 & _T_390; // @[MemPrimitives.scala 110:228:@19006.4]
  assign _T_523 = _T_436 & _T_396; // @[MemPrimitives.scala 110:228:@19010.4]
  assign _T_529 = _T_442 & _T_402; // @[MemPrimitives.scala 110:228:@19014.4]
  assign _T_531 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@19023.4]
  assign _T_532 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@19024.4]
  assign _T_533 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@19025.4]
  assign _T_534 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@19026.4]
  assign _T_536 = {_T_531,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19028.4]
  assign _T_538 = {_T_532,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19030.4]
  assign _T_540 = {_T_533,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19032.4]
  assign _T_542 = {_T_534,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19034.4]
  assign _T_543 = _T_533 ? _T_540 : _T_542; // @[Mux.scala 31:69:@19035.4]
  assign _T_544 = _T_532 ? _T_538 : _T_543; // @[Mux.scala 31:69:@19036.4]
  assign _T_545 = _T_531 ? _T_536 : _T_544; // @[Mux.scala 31:69:@19037.4]
  assign _T_550 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19044.4]
  assign _T_553 = _T_550 & _T_300; // @[MemPrimitives.scala 110:228:@19046.4]
  assign _T_556 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19048.4]
  assign _T_559 = _T_556 & _T_306; // @[MemPrimitives.scala 110:228:@19050.4]
  assign _T_562 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19052.4]
  assign _T_565 = _T_562 & _T_312; // @[MemPrimitives.scala 110:228:@19054.4]
  assign _T_568 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19056.4]
  assign _T_571 = _T_568 & _T_318; // @[MemPrimitives.scala 110:228:@19058.4]
  assign _T_573 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@19067.4]
  assign _T_574 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@19068.4]
  assign _T_575 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@19069.4]
  assign _T_576 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@19070.4]
  assign _T_578 = {_T_573,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19072.4]
  assign _T_580 = {_T_574,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19074.4]
  assign _T_582 = {_T_575,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19076.4]
  assign _T_584 = {_T_576,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19078.4]
  assign _T_585 = _T_575 ? _T_582 : _T_584; // @[Mux.scala 31:69:@19079.4]
  assign _T_586 = _T_574 ? _T_580 : _T_585; // @[Mux.scala 31:69:@19080.4]
  assign _T_587 = _T_573 ? _T_578 : _T_586; // @[Mux.scala 31:69:@19081.4]
  assign _T_595 = _T_550 & _T_342; // @[MemPrimitives.scala 110:228:@19090.4]
  assign _T_601 = _T_556 & _T_348; // @[MemPrimitives.scala 110:228:@19094.4]
  assign _T_607 = _T_562 & _T_354; // @[MemPrimitives.scala 110:228:@19098.4]
  assign _T_613 = _T_568 & _T_360; // @[MemPrimitives.scala 110:228:@19102.4]
  assign _T_615 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@19111.4]
  assign _T_616 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@19112.4]
  assign _T_617 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@19113.4]
  assign _T_618 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@19114.4]
  assign _T_620 = {_T_615,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19116.4]
  assign _T_622 = {_T_616,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19118.4]
  assign _T_624 = {_T_617,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19120.4]
  assign _T_626 = {_T_618,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19122.4]
  assign _T_627 = _T_617 ? _T_624 : _T_626; // @[Mux.scala 31:69:@19123.4]
  assign _T_628 = _T_616 ? _T_622 : _T_627; // @[Mux.scala 31:69:@19124.4]
  assign _T_629 = _T_615 ? _T_620 : _T_628; // @[Mux.scala 31:69:@19125.4]
  assign _T_637 = _T_550 & _T_384; // @[MemPrimitives.scala 110:228:@19134.4]
  assign _T_643 = _T_556 & _T_390; // @[MemPrimitives.scala 110:228:@19138.4]
  assign _T_649 = _T_562 & _T_396; // @[MemPrimitives.scala 110:228:@19142.4]
  assign _T_655 = _T_568 & _T_402; // @[MemPrimitives.scala 110:228:@19146.4]
  assign _T_657 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@19155.4]
  assign _T_658 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@19156.4]
  assign _T_659 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@19157.4]
  assign _T_660 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@19158.4]
  assign _T_662 = {_T_657,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19160.4]
  assign _T_664 = {_T_658,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19162.4]
  assign _T_666 = {_T_659,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19164.4]
  assign _T_668 = {_T_660,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19166.4]
  assign _T_669 = _T_659 ? _T_666 : _T_668; // @[Mux.scala 31:69:@19167.4]
  assign _T_670 = _T_658 ? _T_664 : _T_669; // @[Mux.scala 31:69:@19168.4]
  assign _T_671 = _T_657 ? _T_662 : _T_670; // @[Mux.scala 31:69:@19169.4]
  assign _T_676 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19176.4]
  assign _T_679 = _T_676 & _T_300; // @[MemPrimitives.scala 110:228:@19178.4]
  assign _T_682 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19180.4]
  assign _T_685 = _T_682 & _T_306; // @[MemPrimitives.scala 110:228:@19182.4]
  assign _T_688 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19184.4]
  assign _T_691 = _T_688 & _T_312; // @[MemPrimitives.scala 110:228:@19186.4]
  assign _T_694 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19188.4]
  assign _T_697 = _T_694 & _T_318; // @[MemPrimitives.scala 110:228:@19190.4]
  assign _T_699 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@19199.4]
  assign _T_700 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@19200.4]
  assign _T_701 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@19201.4]
  assign _T_702 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@19202.4]
  assign _T_704 = {_T_699,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19204.4]
  assign _T_706 = {_T_700,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19206.4]
  assign _T_708 = {_T_701,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19208.4]
  assign _T_710 = {_T_702,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19210.4]
  assign _T_711 = _T_701 ? _T_708 : _T_710; // @[Mux.scala 31:69:@19211.4]
  assign _T_712 = _T_700 ? _T_706 : _T_711; // @[Mux.scala 31:69:@19212.4]
  assign _T_713 = _T_699 ? _T_704 : _T_712; // @[Mux.scala 31:69:@19213.4]
  assign _T_721 = _T_676 & _T_342; // @[MemPrimitives.scala 110:228:@19222.4]
  assign _T_727 = _T_682 & _T_348; // @[MemPrimitives.scala 110:228:@19226.4]
  assign _T_733 = _T_688 & _T_354; // @[MemPrimitives.scala 110:228:@19230.4]
  assign _T_739 = _T_694 & _T_360; // @[MemPrimitives.scala 110:228:@19234.4]
  assign _T_741 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@19243.4]
  assign _T_742 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@19244.4]
  assign _T_743 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@19245.4]
  assign _T_744 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@19246.4]
  assign _T_746 = {_T_741,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19248.4]
  assign _T_748 = {_T_742,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19250.4]
  assign _T_750 = {_T_743,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19252.4]
  assign _T_752 = {_T_744,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19254.4]
  assign _T_753 = _T_743 ? _T_750 : _T_752; // @[Mux.scala 31:69:@19255.4]
  assign _T_754 = _T_742 ? _T_748 : _T_753; // @[Mux.scala 31:69:@19256.4]
  assign _T_755 = _T_741 ? _T_746 : _T_754; // @[Mux.scala 31:69:@19257.4]
  assign _T_763 = _T_676 & _T_384; // @[MemPrimitives.scala 110:228:@19266.4]
  assign _T_769 = _T_682 & _T_390; // @[MemPrimitives.scala 110:228:@19270.4]
  assign _T_775 = _T_688 & _T_396; // @[MemPrimitives.scala 110:228:@19274.4]
  assign _T_781 = _T_694 & _T_402; // @[MemPrimitives.scala 110:228:@19278.4]
  assign _T_783 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@19287.4]
  assign _T_784 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@19288.4]
  assign _T_785 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@19289.4]
  assign _T_786 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@19290.4]
  assign _T_788 = {_T_783,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19292.4]
  assign _T_790 = {_T_784,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19294.4]
  assign _T_792 = {_T_785,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19296.4]
  assign _T_794 = {_T_786,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19298.4]
  assign _T_795 = _T_785 ? _T_792 : _T_794; // @[Mux.scala 31:69:@19299.4]
  assign _T_796 = _T_784 ? _T_790 : _T_795; // @[Mux.scala 31:69:@19300.4]
  assign _T_797 = _T_783 ? _T_788 : _T_796; // @[Mux.scala 31:69:@19301.4]
  assign _T_893 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@19430.4 package.scala 96:25:@19431.4]
  assign _T_897 = _T_893 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19440.4]
  assign _T_890 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@19422.4 package.scala 96:25:@19423.4]
  assign _T_898 = _T_890 ? Mem1D_9_io_output : _T_897; // @[Mux.scala 31:69:@19441.4]
  assign _T_887 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@19414.4 package.scala 96:25:@19415.4]
  assign _T_899 = _T_887 ? Mem1D_8_io_output : _T_898; // @[Mux.scala 31:69:@19442.4]
  assign _T_884 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@19406.4 package.scala 96:25:@19407.4]
  assign _T_900 = _T_884 ? Mem1D_7_io_output : _T_899; // @[Mux.scala 31:69:@19443.4]
  assign _T_881 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@19398.4 package.scala 96:25:@19399.4]
  assign _T_901 = _T_881 ? Mem1D_6_io_output : _T_900; // @[Mux.scala 31:69:@19444.4]
  assign _T_878 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@19390.4 package.scala 96:25:@19391.4]
  assign _T_902 = _T_878 ? Mem1D_5_io_output : _T_901; // @[Mux.scala 31:69:@19445.4]
  assign _T_875 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@19382.4 package.scala 96:25:@19383.4]
  assign _T_903 = _T_875 ? Mem1D_4_io_output : _T_902; // @[Mux.scala 31:69:@19446.4]
  assign _T_872 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@19374.4 package.scala 96:25:@19375.4]
  assign _T_904 = _T_872 ? Mem1D_3_io_output : _T_903; // @[Mux.scala 31:69:@19447.4]
  assign _T_869 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@19366.4 package.scala 96:25:@19367.4]
  assign _T_905 = _T_869 ? Mem1D_2_io_output : _T_904; // @[Mux.scala 31:69:@19448.4]
  assign _T_866 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@19358.4 package.scala 96:25:@19359.4]
  assign _T_906 = _T_866 ? Mem1D_1_io_output : _T_905; // @[Mux.scala 31:69:@19449.4]
  assign _T_863 = RetimeWrapper_io_out; // @[package.scala 96:25:@19350.4 package.scala 96:25:@19351.4]
  assign _T_1000 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@19574.4 package.scala 96:25:@19575.4]
  assign _T_1004 = _T_1000 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19584.4]
  assign _T_997 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@19566.4 package.scala 96:25:@19567.4]
  assign _T_1005 = _T_997 ? Mem1D_9_io_output : _T_1004; // @[Mux.scala 31:69:@19585.4]
  assign _T_994 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@19558.4 package.scala 96:25:@19559.4]
  assign _T_1006 = _T_994 ? Mem1D_8_io_output : _T_1005; // @[Mux.scala 31:69:@19586.4]
  assign _T_991 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@19550.4 package.scala 96:25:@19551.4]
  assign _T_1007 = _T_991 ? Mem1D_7_io_output : _T_1006; // @[Mux.scala 31:69:@19587.4]
  assign _T_988 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@19542.4 package.scala 96:25:@19543.4]
  assign _T_1008 = _T_988 ? Mem1D_6_io_output : _T_1007; // @[Mux.scala 31:69:@19588.4]
  assign _T_985 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@19534.4 package.scala 96:25:@19535.4]
  assign _T_1009 = _T_985 ? Mem1D_5_io_output : _T_1008; // @[Mux.scala 31:69:@19589.4]
  assign _T_982 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@19526.4 package.scala 96:25:@19527.4]
  assign _T_1010 = _T_982 ? Mem1D_4_io_output : _T_1009; // @[Mux.scala 31:69:@19590.4]
  assign _T_979 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@19518.4 package.scala 96:25:@19519.4]
  assign _T_1011 = _T_979 ? Mem1D_3_io_output : _T_1010; // @[Mux.scala 31:69:@19591.4]
  assign _T_976 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@19510.4 package.scala 96:25:@19511.4]
  assign _T_1012 = _T_976 ? Mem1D_2_io_output : _T_1011; // @[Mux.scala 31:69:@19592.4]
  assign _T_973 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@19502.4 package.scala 96:25:@19503.4]
  assign _T_1013 = _T_973 ? Mem1D_1_io_output : _T_1012; // @[Mux.scala 31:69:@19593.4]
  assign _T_970 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@19494.4 package.scala 96:25:@19495.4]
  assign _T_1107 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@19718.4 package.scala 96:25:@19719.4]
  assign _T_1111 = _T_1107 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19728.4]
  assign _T_1104 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@19710.4 package.scala 96:25:@19711.4]
  assign _T_1112 = _T_1104 ? Mem1D_9_io_output : _T_1111; // @[Mux.scala 31:69:@19729.4]
  assign _T_1101 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@19702.4 package.scala 96:25:@19703.4]
  assign _T_1113 = _T_1101 ? Mem1D_8_io_output : _T_1112; // @[Mux.scala 31:69:@19730.4]
  assign _T_1098 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@19694.4 package.scala 96:25:@19695.4]
  assign _T_1114 = _T_1098 ? Mem1D_7_io_output : _T_1113; // @[Mux.scala 31:69:@19731.4]
  assign _T_1095 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@19686.4 package.scala 96:25:@19687.4]
  assign _T_1115 = _T_1095 ? Mem1D_6_io_output : _T_1114; // @[Mux.scala 31:69:@19732.4]
  assign _T_1092 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@19678.4 package.scala 96:25:@19679.4]
  assign _T_1116 = _T_1092 ? Mem1D_5_io_output : _T_1115; // @[Mux.scala 31:69:@19733.4]
  assign _T_1089 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@19670.4 package.scala 96:25:@19671.4]
  assign _T_1117 = _T_1089 ? Mem1D_4_io_output : _T_1116; // @[Mux.scala 31:69:@19734.4]
  assign _T_1086 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@19662.4 package.scala 96:25:@19663.4]
  assign _T_1118 = _T_1086 ? Mem1D_3_io_output : _T_1117; // @[Mux.scala 31:69:@19735.4]
  assign _T_1083 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@19654.4 package.scala 96:25:@19655.4]
  assign _T_1119 = _T_1083 ? Mem1D_2_io_output : _T_1118; // @[Mux.scala 31:69:@19736.4]
  assign _T_1080 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@19646.4 package.scala 96:25:@19647.4]
  assign _T_1120 = _T_1080 ? Mem1D_1_io_output : _T_1119; // @[Mux.scala 31:69:@19737.4]
  assign _T_1077 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@19638.4 package.scala 96:25:@19639.4]
  assign _T_1214 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@19862.4 package.scala 96:25:@19863.4]
  assign _T_1218 = _T_1214 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@19872.4]
  assign _T_1211 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@19854.4 package.scala 96:25:@19855.4]
  assign _T_1219 = _T_1211 ? Mem1D_9_io_output : _T_1218; // @[Mux.scala 31:69:@19873.4]
  assign _T_1208 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@19846.4 package.scala 96:25:@19847.4]
  assign _T_1220 = _T_1208 ? Mem1D_8_io_output : _T_1219; // @[Mux.scala 31:69:@19874.4]
  assign _T_1205 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@19838.4 package.scala 96:25:@19839.4]
  assign _T_1221 = _T_1205 ? Mem1D_7_io_output : _T_1220; // @[Mux.scala 31:69:@19875.4]
  assign _T_1202 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@19830.4 package.scala 96:25:@19831.4]
  assign _T_1222 = _T_1202 ? Mem1D_6_io_output : _T_1221; // @[Mux.scala 31:69:@19876.4]
  assign _T_1199 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@19822.4 package.scala 96:25:@19823.4]
  assign _T_1223 = _T_1199 ? Mem1D_5_io_output : _T_1222; // @[Mux.scala 31:69:@19877.4]
  assign _T_1196 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@19814.4 package.scala 96:25:@19815.4]
  assign _T_1224 = _T_1196 ? Mem1D_4_io_output : _T_1223; // @[Mux.scala 31:69:@19878.4]
  assign _T_1193 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@19806.4 package.scala 96:25:@19807.4]
  assign _T_1225 = _T_1193 ? Mem1D_3_io_output : _T_1224; // @[Mux.scala 31:69:@19879.4]
  assign _T_1190 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@19798.4 package.scala 96:25:@19799.4]
  assign _T_1226 = _T_1190 ? Mem1D_2_io_output : _T_1225; // @[Mux.scala 31:69:@19880.4]
  assign _T_1187 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@19790.4 package.scala 96:25:@19791.4]
  assign _T_1227 = _T_1187 ? Mem1D_1_io_output : _T_1226; // @[Mux.scala 31:69:@19881.4]
  assign _T_1184 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@19782.4 package.scala 96:25:@19783.4]
  assign io_rPort_3_output_0 = _T_1184 ? Mem1D_io_output : _T_1227; // @[MemPrimitives.scala 152:13:@19883.4]
  assign io_rPort_2_output_0 = _T_1077 ? Mem1D_io_output : _T_1120; // @[MemPrimitives.scala 152:13:@19739.4]
  assign io_rPort_1_output_0 = _T_970 ? Mem1D_io_output : _T_1013; // @[MemPrimitives.scala 152:13:@19595.4]
  assign io_rPort_0_output_0 = _T_863 ? Mem1D_io_output : _T_906; // @[MemPrimitives.scala 152:13:@19451.4]
  assign Mem1D_clock = clock; // @[:@18445.4]
  assign Mem1D_reset = reset; // @[:@18446.4]
  assign Mem1D_io_r_ofs_0 = _T_335[9:0]; // @[MemPrimitives.scala 131:28:@18821.4]
  assign Mem1D_io_r_backpressure = _T_335[10]; // @[MemPrimitives.scala 132:32:@18822.4]
  assign Mem1D_io_w_ofs_0 = _T_172[9:0]; // @[MemPrimitives.scala 94:28:@18645.4]
  assign Mem1D_io_w_data_0 = _T_172[41:10]; // @[MemPrimitives.scala 95:29:@18646.4]
  assign Mem1D_io_w_en_0 = _T_172[42]; // @[MemPrimitives.scala 96:27:@18647.4]
  assign Mem1D_1_clock = clock; // @[:@18461.4]
  assign Mem1D_1_reset = reset; // @[:@18462.4]
  assign Mem1D_1_io_r_ofs_0 = _T_377[9:0]; // @[MemPrimitives.scala 131:28:@18865.4]
  assign Mem1D_1_io_r_backpressure = _T_377[10]; // @[MemPrimitives.scala 132:32:@18866.4]
  assign Mem1D_1_io_w_ofs_0 = _T_183[9:0]; // @[MemPrimitives.scala 94:28:@18657.4]
  assign Mem1D_1_io_w_data_0 = _T_183[41:10]; // @[MemPrimitives.scala 95:29:@18658.4]
  assign Mem1D_1_io_w_en_0 = _T_183[42]; // @[MemPrimitives.scala 96:27:@18659.4]
  assign Mem1D_2_clock = clock; // @[:@18477.4]
  assign Mem1D_2_reset = reset; // @[:@18478.4]
  assign Mem1D_2_io_r_ofs_0 = _T_419[9:0]; // @[MemPrimitives.scala 131:28:@18909.4]
  assign Mem1D_2_io_r_backpressure = _T_419[10]; // @[MemPrimitives.scala 132:32:@18910.4]
  assign Mem1D_2_io_w_ofs_0 = _T_194[9:0]; // @[MemPrimitives.scala 94:28:@18669.4]
  assign Mem1D_2_io_w_data_0 = _T_194[41:10]; // @[MemPrimitives.scala 95:29:@18670.4]
  assign Mem1D_2_io_w_en_0 = _T_194[42]; // @[MemPrimitives.scala 96:27:@18671.4]
  assign Mem1D_3_clock = clock; // @[:@18493.4]
  assign Mem1D_3_reset = reset; // @[:@18494.4]
  assign Mem1D_3_io_r_ofs_0 = _T_461[9:0]; // @[MemPrimitives.scala 131:28:@18953.4]
  assign Mem1D_3_io_r_backpressure = _T_461[10]; // @[MemPrimitives.scala 132:32:@18954.4]
  assign Mem1D_3_io_w_ofs_0 = _T_205[9:0]; // @[MemPrimitives.scala 94:28:@18681.4]
  assign Mem1D_3_io_w_data_0 = _T_205[41:10]; // @[MemPrimitives.scala 95:29:@18682.4]
  assign Mem1D_3_io_w_en_0 = _T_205[42]; // @[MemPrimitives.scala 96:27:@18683.4]
  assign Mem1D_4_clock = clock; // @[:@18509.4]
  assign Mem1D_4_reset = reset; // @[:@18510.4]
  assign Mem1D_4_io_r_ofs_0 = _T_503[9:0]; // @[MemPrimitives.scala 131:28:@18997.4]
  assign Mem1D_4_io_r_backpressure = _T_503[10]; // @[MemPrimitives.scala 132:32:@18998.4]
  assign Mem1D_4_io_w_ofs_0 = _T_216[9:0]; // @[MemPrimitives.scala 94:28:@18693.4]
  assign Mem1D_4_io_w_data_0 = _T_216[41:10]; // @[MemPrimitives.scala 95:29:@18694.4]
  assign Mem1D_4_io_w_en_0 = _T_216[42]; // @[MemPrimitives.scala 96:27:@18695.4]
  assign Mem1D_5_clock = clock; // @[:@18525.4]
  assign Mem1D_5_reset = reset; // @[:@18526.4]
  assign Mem1D_5_io_r_ofs_0 = _T_545[9:0]; // @[MemPrimitives.scala 131:28:@19041.4]
  assign Mem1D_5_io_r_backpressure = _T_545[10]; // @[MemPrimitives.scala 132:32:@19042.4]
  assign Mem1D_5_io_w_ofs_0 = _T_227[9:0]; // @[MemPrimitives.scala 94:28:@18705.4]
  assign Mem1D_5_io_w_data_0 = _T_227[41:10]; // @[MemPrimitives.scala 95:29:@18706.4]
  assign Mem1D_5_io_w_en_0 = _T_227[42]; // @[MemPrimitives.scala 96:27:@18707.4]
  assign Mem1D_6_clock = clock; // @[:@18541.4]
  assign Mem1D_6_reset = reset; // @[:@18542.4]
  assign Mem1D_6_io_r_ofs_0 = _T_587[9:0]; // @[MemPrimitives.scala 131:28:@19085.4]
  assign Mem1D_6_io_r_backpressure = _T_587[10]; // @[MemPrimitives.scala 132:32:@19086.4]
  assign Mem1D_6_io_w_ofs_0 = _T_238[9:0]; // @[MemPrimitives.scala 94:28:@18717.4]
  assign Mem1D_6_io_w_data_0 = _T_238[41:10]; // @[MemPrimitives.scala 95:29:@18718.4]
  assign Mem1D_6_io_w_en_0 = _T_238[42]; // @[MemPrimitives.scala 96:27:@18719.4]
  assign Mem1D_7_clock = clock; // @[:@18557.4]
  assign Mem1D_7_reset = reset; // @[:@18558.4]
  assign Mem1D_7_io_r_ofs_0 = _T_629[9:0]; // @[MemPrimitives.scala 131:28:@19129.4]
  assign Mem1D_7_io_r_backpressure = _T_629[10]; // @[MemPrimitives.scala 132:32:@19130.4]
  assign Mem1D_7_io_w_ofs_0 = _T_249[9:0]; // @[MemPrimitives.scala 94:28:@18729.4]
  assign Mem1D_7_io_w_data_0 = _T_249[41:10]; // @[MemPrimitives.scala 95:29:@18730.4]
  assign Mem1D_7_io_w_en_0 = _T_249[42]; // @[MemPrimitives.scala 96:27:@18731.4]
  assign Mem1D_8_clock = clock; // @[:@18573.4]
  assign Mem1D_8_reset = reset; // @[:@18574.4]
  assign Mem1D_8_io_r_ofs_0 = _T_671[9:0]; // @[MemPrimitives.scala 131:28:@19173.4]
  assign Mem1D_8_io_r_backpressure = _T_671[10]; // @[MemPrimitives.scala 132:32:@19174.4]
  assign Mem1D_8_io_w_ofs_0 = _T_260[9:0]; // @[MemPrimitives.scala 94:28:@18741.4]
  assign Mem1D_8_io_w_data_0 = _T_260[41:10]; // @[MemPrimitives.scala 95:29:@18742.4]
  assign Mem1D_8_io_w_en_0 = _T_260[42]; // @[MemPrimitives.scala 96:27:@18743.4]
  assign Mem1D_9_clock = clock; // @[:@18589.4]
  assign Mem1D_9_reset = reset; // @[:@18590.4]
  assign Mem1D_9_io_r_ofs_0 = _T_713[9:0]; // @[MemPrimitives.scala 131:28:@19217.4]
  assign Mem1D_9_io_r_backpressure = _T_713[10]; // @[MemPrimitives.scala 132:32:@19218.4]
  assign Mem1D_9_io_w_ofs_0 = _T_271[9:0]; // @[MemPrimitives.scala 94:28:@18753.4]
  assign Mem1D_9_io_w_data_0 = _T_271[41:10]; // @[MemPrimitives.scala 95:29:@18754.4]
  assign Mem1D_9_io_w_en_0 = _T_271[42]; // @[MemPrimitives.scala 96:27:@18755.4]
  assign Mem1D_10_clock = clock; // @[:@18605.4]
  assign Mem1D_10_reset = reset; // @[:@18606.4]
  assign Mem1D_10_io_r_ofs_0 = _T_755[9:0]; // @[MemPrimitives.scala 131:28:@19261.4]
  assign Mem1D_10_io_r_backpressure = _T_755[10]; // @[MemPrimitives.scala 132:32:@19262.4]
  assign Mem1D_10_io_w_ofs_0 = _T_282[9:0]; // @[MemPrimitives.scala 94:28:@18765.4]
  assign Mem1D_10_io_w_data_0 = _T_282[41:10]; // @[MemPrimitives.scala 95:29:@18766.4]
  assign Mem1D_10_io_w_en_0 = _T_282[42]; // @[MemPrimitives.scala 96:27:@18767.4]
  assign Mem1D_11_clock = clock; // @[:@18621.4]
  assign Mem1D_11_reset = reset; // @[:@18622.4]
  assign Mem1D_11_io_r_ofs_0 = _T_797[9:0]; // @[MemPrimitives.scala 131:28:@19305.4]
  assign Mem1D_11_io_r_backpressure = _T_797[10]; // @[MemPrimitives.scala 132:32:@19306.4]
  assign Mem1D_11_io_w_ofs_0 = _T_293[9:0]; // @[MemPrimitives.scala 94:28:@18777.4]
  assign Mem1D_11_io_w_data_0 = _T_293[41:10]; // @[MemPrimitives.scala 95:29:@18778.4]
  assign Mem1D_11_io_w_en_0 = _T_293[42]; // @[MemPrimitives.scala 96:27:@18779.4]
  assign StickySelects_clock = clock; // @[:@18797.4]
  assign StickySelects_reset = reset; // @[:@18798.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_301; // @[MemPrimitives.scala 125:64:@18799.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_307; // @[MemPrimitives.scala 125:64:@18800.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_313; // @[MemPrimitives.scala 125:64:@18801.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_319; // @[MemPrimitives.scala 125:64:@18802.4]
  assign StickySelects_1_clock = clock; // @[:@18841.4]
  assign StickySelects_1_reset = reset; // @[:@18842.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_343; // @[MemPrimitives.scala 125:64:@18843.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_349; // @[MemPrimitives.scala 125:64:@18844.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_355; // @[MemPrimitives.scala 125:64:@18845.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_361; // @[MemPrimitives.scala 125:64:@18846.4]
  assign StickySelects_2_clock = clock; // @[:@18885.4]
  assign StickySelects_2_reset = reset; // @[:@18886.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_385; // @[MemPrimitives.scala 125:64:@18887.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_391; // @[MemPrimitives.scala 125:64:@18888.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_397; // @[MemPrimitives.scala 125:64:@18889.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_403; // @[MemPrimitives.scala 125:64:@18890.4]
  assign StickySelects_3_clock = clock; // @[:@18929.4]
  assign StickySelects_3_reset = reset; // @[:@18930.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_427; // @[MemPrimitives.scala 125:64:@18931.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_433; // @[MemPrimitives.scala 125:64:@18932.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_439; // @[MemPrimitives.scala 125:64:@18933.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_445; // @[MemPrimitives.scala 125:64:@18934.4]
  assign StickySelects_4_clock = clock; // @[:@18973.4]
  assign StickySelects_4_reset = reset; // @[:@18974.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_469; // @[MemPrimitives.scala 125:64:@18975.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_475; // @[MemPrimitives.scala 125:64:@18976.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_481; // @[MemPrimitives.scala 125:64:@18977.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_487; // @[MemPrimitives.scala 125:64:@18978.4]
  assign StickySelects_5_clock = clock; // @[:@19017.4]
  assign StickySelects_5_reset = reset; // @[:@19018.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_511; // @[MemPrimitives.scala 125:64:@19019.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_517; // @[MemPrimitives.scala 125:64:@19020.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_523; // @[MemPrimitives.scala 125:64:@19021.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_529; // @[MemPrimitives.scala 125:64:@19022.4]
  assign StickySelects_6_clock = clock; // @[:@19061.4]
  assign StickySelects_6_reset = reset; // @[:@19062.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_553; // @[MemPrimitives.scala 125:64:@19063.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_559; // @[MemPrimitives.scala 125:64:@19064.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_565; // @[MemPrimitives.scala 125:64:@19065.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_571; // @[MemPrimitives.scala 125:64:@19066.4]
  assign StickySelects_7_clock = clock; // @[:@19105.4]
  assign StickySelects_7_reset = reset; // @[:@19106.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_595; // @[MemPrimitives.scala 125:64:@19107.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_601; // @[MemPrimitives.scala 125:64:@19108.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_607; // @[MemPrimitives.scala 125:64:@19109.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_613; // @[MemPrimitives.scala 125:64:@19110.4]
  assign StickySelects_8_clock = clock; // @[:@19149.4]
  assign StickySelects_8_reset = reset; // @[:@19150.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_637; // @[MemPrimitives.scala 125:64:@19151.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_643; // @[MemPrimitives.scala 125:64:@19152.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_649; // @[MemPrimitives.scala 125:64:@19153.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_655; // @[MemPrimitives.scala 125:64:@19154.4]
  assign StickySelects_9_clock = clock; // @[:@19193.4]
  assign StickySelects_9_reset = reset; // @[:@19194.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_679; // @[MemPrimitives.scala 125:64:@19195.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 125:64:@19196.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_691; // @[MemPrimitives.scala 125:64:@19197.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_697; // @[MemPrimitives.scala 125:64:@19198.4]
  assign StickySelects_10_clock = clock; // @[:@19237.4]
  assign StickySelects_10_reset = reset; // @[:@19238.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_721; // @[MemPrimitives.scala 125:64:@19239.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@19240.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@19241.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@19242.4]
  assign StickySelects_11_clock = clock; // @[:@19281.4]
  assign StickySelects_11_reset = reset; // @[:@19282.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@19283.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@19284.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_775; // @[MemPrimitives.scala 125:64:@19285.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_781; // @[MemPrimitives.scala 125:64:@19286.4]
  assign RetimeWrapper_clock = clock; // @[:@19346.4]
  assign RetimeWrapper_reset = reset; // @[:@19347.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19349.4]
  assign RetimeWrapper_io_in = _T_301 & io_rPort_0_en_0; // @[package.scala 94:16:@19348.4]
  assign RetimeWrapper_1_clock = clock; // @[:@19354.4]
  assign RetimeWrapper_1_reset = reset; // @[:@19355.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19357.4]
  assign RetimeWrapper_1_io_in = _T_343 & io_rPort_0_en_0; // @[package.scala 94:16:@19356.4]
  assign RetimeWrapper_2_clock = clock; // @[:@19362.4]
  assign RetimeWrapper_2_reset = reset; // @[:@19363.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19365.4]
  assign RetimeWrapper_2_io_in = _T_385 & io_rPort_0_en_0; // @[package.scala 94:16:@19364.4]
  assign RetimeWrapper_3_clock = clock; // @[:@19370.4]
  assign RetimeWrapper_3_reset = reset; // @[:@19371.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19373.4]
  assign RetimeWrapper_3_io_in = _T_427 & io_rPort_0_en_0; // @[package.scala 94:16:@19372.4]
  assign RetimeWrapper_4_clock = clock; // @[:@19378.4]
  assign RetimeWrapper_4_reset = reset; // @[:@19379.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19381.4]
  assign RetimeWrapper_4_io_in = _T_469 & io_rPort_0_en_0; // @[package.scala 94:16:@19380.4]
  assign RetimeWrapper_5_clock = clock; // @[:@19386.4]
  assign RetimeWrapper_5_reset = reset; // @[:@19387.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19389.4]
  assign RetimeWrapper_5_io_in = _T_511 & io_rPort_0_en_0; // @[package.scala 94:16:@19388.4]
  assign RetimeWrapper_6_clock = clock; // @[:@19394.4]
  assign RetimeWrapper_6_reset = reset; // @[:@19395.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19397.4]
  assign RetimeWrapper_6_io_in = _T_553 & io_rPort_0_en_0; // @[package.scala 94:16:@19396.4]
  assign RetimeWrapper_7_clock = clock; // @[:@19402.4]
  assign RetimeWrapper_7_reset = reset; // @[:@19403.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19405.4]
  assign RetimeWrapper_7_io_in = _T_595 & io_rPort_0_en_0; // @[package.scala 94:16:@19404.4]
  assign RetimeWrapper_8_clock = clock; // @[:@19410.4]
  assign RetimeWrapper_8_reset = reset; // @[:@19411.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19413.4]
  assign RetimeWrapper_8_io_in = _T_637 & io_rPort_0_en_0; // @[package.scala 94:16:@19412.4]
  assign RetimeWrapper_9_clock = clock; // @[:@19418.4]
  assign RetimeWrapper_9_reset = reset; // @[:@19419.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19421.4]
  assign RetimeWrapper_9_io_in = _T_679 & io_rPort_0_en_0; // @[package.scala 94:16:@19420.4]
  assign RetimeWrapper_10_clock = clock; // @[:@19426.4]
  assign RetimeWrapper_10_reset = reset; // @[:@19427.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19429.4]
  assign RetimeWrapper_10_io_in = _T_721 & io_rPort_0_en_0; // @[package.scala 94:16:@19428.4]
  assign RetimeWrapper_11_clock = clock; // @[:@19434.4]
  assign RetimeWrapper_11_reset = reset; // @[:@19435.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19437.4]
  assign RetimeWrapper_11_io_in = _T_763 & io_rPort_0_en_0; // @[package.scala 94:16:@19436.4]
  assign RetimeWrapper_12_clock = clock; // @[:@19490.4]
  assign RetimeWrapper_12_reset = reset; // @[:@19491.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19493.4]
  assign RetimeWrapper_12_io_in = _T_307 & io_rPort_1_en_0; // @[package.scala 94:16:@19492.4]
  assign RetimeWrapper_13_clock = clock; // @[:@19498.4]
  assign RetimeWrapper_13_reset = reset; // @[:@19499.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19501.4]
  assign RetimeWrapper_13_io_in = _T_349 & io_rPort_1_en_0; // @[package.scala 94:16:@19500.4]
  assign RetimeWrapper_14_clock = clock; // @[:@19506.4]
  assign RetimeWrapper_14_reset = reset; // @[:@19507.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19509.4]
  assign RetimeWrapper_14_io_in = _T_391 & io_rPort_1_en_0; // @[package.scala 94:16:@19508.4]
  assign RetimeWrapper_15_clock = clock; // @[:@19514.4]
  assign RetimeWrapper_15_reset = reset; // @[:@19515.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19517.4]
  assign RetimeWrapper_15_io_in = _T_433 & io_rPort_1_en_0; // @[package.scala 94:16:@19516.4]
  assign RetimeWrapper_16_clock = clock; // @[:@19522.4]
  assign RetimeWrapper_16_reset = reset; // @[:@19523.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19525.4]
  assign RetimeWrapper_16_io_in = _T_475 & io_rPort_1_en_0; // @[package.scala 94:16:@19524.4]
  assign RetimeWrapper_17_clock = clock; // @[:@19530.4]
  assign RetimeWrapper_17_reset = reset; // @[:@19531.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19533.4]
  assign RetimeWrapper_17_io_in = _T_517 & io_rPort_1_en_0; // @[package.scala 94:16:@19532.4]
  assign RetimeWrapper_18_clock = clock; // @[:@19538.4]
  assign RetimeWrapper_18_reset = reset; // @[:@19539.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19541.4]
  assign RetimeWrapper_18_io_in = _T_559 & io_rPort_1_en_0; // @[package.scala 94:16:@19540.4]
  assign RetimeWrapper_19_clock = clock; // @[:@19546.4]
  assign RetimeWrapper_19_reset = reset; // @[:@19547.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19549.4]
  assign RetimeWrapper_19_io_in = _T_601 & io_rPort_1_en_0; // @[package.scala 94:16:@19548.4]
  assign RetimeWrapper_20_clock = clock; // @[:@19554.4]
  assign RetimeWrapper_20_reset = reset; // @[:@19555.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19557.4]
  assign RetimeWrapper_20_io_in = _T_643 & io_rPort_1_en_0; // @[package.scala 94:16:@19556.4]
  assign RetimeWrapper_21_clock = clock; // @[:@19562.4]
  assign RetimeWrapper_21_reset = reset; // @[:@19563.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19565.4]
  assign RetimeWrapper_21_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@19564.4]
  assign RetimeWrapper_22_clock = clock; // @[:@19570.4]
  assign RetimeWrapper_22_reset = reset; // @[:@19571.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19573.4]
  assign RetimeWrapper_22_io_in = _T_727 & io_rPort_1_en_0; // @[package.scala 94:16:@19572.4]
  assign RetimeWrapper_23_clock = clock; // @[:@19578.4]
  assign RetimeWrapper_23_reset = reset; // @[:@19579.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19581.4]
  assign RetimeWrapper_23_io_in = _T_769 & io_rPort_1_en_0; // @[package.scala 94:16:@19580.4]
  assign RetimeWrapper_24_clock = clock; // @[:@19634.4]
  assign RetimeWrapper_24_reset = reset; // @[:@19635.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19637.4]
  assign RetimeWrapper_24_io_in = _T_313 & io_rPort_2_en_0; // @[package.scala 94:16:@19636.4]
  assign RetimeWrapper_25_clock = clock; // @[:@19642.4]
  assign RetimeWrapper_25_reset = reset; // @[:@19643.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19645.4]
  assign RetimeWrapper_25_io_in = _T_355 & io_rPort_2_en_0; // @[package.scala 94:16:@19644.4]
  assign RetimeWrapper_26_clock = clock; // @[:@19650.4]
  assign RetimeWrapper_26_reset = reset; // @[:@19651.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19653.4]
  assign RetimeWrapper_26_io_in = _T_397 & io_rPort_2_en_0; // @[package.scala 94:16:@19652.4]
  assign RetimeWrapper_27_clock = clock; // @[:@19658.4]
  assign RetimeWrapper_27_reset = reset; // @[:@19659.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19661.4]
  assign RetimeWrapper_27_io_in = _T_439 & io_rPort_2_en_0; // @[package.scala 94:16:@19660.4]
  assign RetimeWrapper_28_clock = clock; // @[:@19666.4]
  assign RetimeWrapper_28_reset = reset; // @[:@19667.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19669.4]
  assign RetimeWrapper_28_io_in = _T_481 & io_rPort_2_en_0; // @[package.scala 94:16:@19668.4]
  assign RetimeWrapper_29_clock = clock; // @[:@19674.4]
  assign RetimeWrapper_29_reset = reset; // @[:@19675.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19677.4]
  assign RetimeWrapper_29_io_in = _T_523 & io_rPort_2_en_0; // @[package.scala 94:16:@19676.4]
  assign RetimeWrapper_30_clock = clock; // @[:@19682.4]
  assign RetimeWrapper_30_reset = reset; // @[:@19683.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19685.4]
  assign RetimeWrapper_30_io_in = _T_565 & io_rPort_2_en_0; // @[package.scala 94:16:@19684.4]
  assign RetimeWrapper_31_clock = clock; // @[:@19690.4]
  assign RetimeWrapper_31_reset = reset; // @[:@19691.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19693.4]
  assign RetimeWrapper_31_io_in = _T_607 & io_rPort_2_en_0; // @[package.scala 94:16:@19692.4]
  assign RetimeWrapper_32_clock = clock; // @[:@19698.4]
  assign RetimeWrapper_32_reset = reset; // @[:@19699.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19701.4]
  assign RetimeWrapper_32_io_in = _T_649 & io_rPort_2_en_0; // @[package.scala 94:16:@19700.4]
  assign RetimeWrapper_33_clock = clock; // @[:@19706.4]
  assign RetimeWrapper_33_reset = reset; // @[:@19707.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19709.4]
  assign RetimeWrapper_33_io_in = _T_691 & io_rPort_2_en_0; // @[package.scala 94:16:@19708.4]
  assign RetimeWrapper_34_clock = clock; // @[:@19714.4]
  assign RetimeWrapper_34_reset = reset; // @[:@19715.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19717.4]
  assign RetimeWrapper_34_io_in = _T_733 & io_rPort_2_en_0; // @[package.scala 94:16:@19716.4]
  assign RetimeWrapper_35_clock = clock; // @[:@19722.4]
  assign RetimeWrapper_35_reset = reset; // @[:@19723.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19725.4]
  assign RetimeWrapper_35_io_in = _T_775 & io_rPort_2_en_0; // @[package.scala 94:16:@19724.4]
  assign RetimeWrapper_36_clock = clock; // @[:@19778.4]
  assign RetimeWrapper_36_reset = reset; // @[:@19779.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19781.4]
  assign RetimeWrapper_36_io_in = _T_319 & io_rPort_3_en_0; // @[package.scala 94:16:@19780.4]
  assign RetimeWrapper_37_clock = clock; // @[:@19786.4]
  assign RetimeWrapper_37_reset = reset; // @[:@19787.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19789.4]
  assign RetimeWrapper_37_io_in = _T_361 & io_rPort_3_en_0; // @[package.scala 94:16:@19788.4]
  assign RetimeWrapper_38_clock = clock; // @[:@19794.4]
  assign RetimeWrapper_38_reset = reset; // @[:@19795.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19797.4]
  assign RetimeWrapper_38_io_in = _T_403 & io_rPort_3_en_0; // @[package.scala 94:16:@19796.4]
  assign RetimeWrapper_39_clock = clock; // @[:@19802.4]
  assign RetimeWrapper_39_reset = reset; // @[:@19803.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19805.4]
  assign RetimeWrapper_39_io_in = _T_445 & io_rPort_3_en_0; // @[package.scala 94:16:@19804.4]
  assign RetimeWrapper_40_clock = clock; // @[:@19810.4]
  assign RetimeWrapper_40_reset = reset; // @[:@19811.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19813.4]
  assign RetimeWrapper_40_io_in = _T_487 & io_rPort_3_en_0; // @[package.scala 94:16:@19812.4]
  assign RetimeWrapper_41_clock = clock; // @[:@19818.4]
  assign RetimeWrapper_41_reset = reset; // @[:@19819.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19821.4]
  assign RetimeWrapper_41_io_in = _T_529 & io_rPort_3_en_0; // @[package.scala 94:16:@19820.4]
  assign RetimeWrapper_42_clock = clock; // @[:@19826.4]
  assign RetimeWrapper_42_reset = reset; // @[:@19827.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19829.4]
  assign RetimeWrapper_42_io_in = _T_571 & io_rPort_3_en_0; // @[package.scala 94:16:@19828.4]
  assign RetimeWrapper_43_clock = clock; // @[:@19834.4]
  assign RetimeWrapper_43_reset = reset; // @[:@19835.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19837.4]
  assign RetimeWrapper_43_io_in = _T_613 & io_rPort_3_en_0; // @[package.scala 94:16:@19836.4]
  assign RetimeWrapper_44_clock = clock; // @[:@19842.4]
  assign RetimeWrapper_44_reset = reset; // @[:@19843.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19845.4]
  assign RetimeWrapper_44_io_in = _T_655 & io_rPort_3_en_0; // @[package.scala 94:16:@19844.4]
  assign RetimeWrapper_45_clock = clock; // @[:@19850.4]
  assign RetimeWrapper_45_reset = reset; // @[:@19851.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19853.4]
  assign RetimeWrapper_45_io_in = _T_697 & io_rPort_3_en_0; // @[package.scala 94:16:@19852.4]
  assign RetimeWrapper_46_clock = clock; // @[:@19858.4]
  assign RetimeWrapper_46_reset = reset; // @[:@19859.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19861.4]
  assign RetimeWrapper_46_io_in = _T_739 & io_rPort_3_en_0; // @[package.scala 94:16:@19860.4]
  assign RetimeWrapper_47_clock = clock; // @[:@19866.4]
  assign RetimeWrapper_47_reset = reset; // @[:@19867.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@19869.4]
  assign RetimeWrapper_47_io_in = _T_781 & io_rPort_3_en_0; // @[package.scala 94:16:@19868.4]
endmodule
module Divider( // @[:@21491.2]
  input         clock, // @[:@21492.4]
  input         io_flow, // @[:@21494.4]
  input  [31:0] io_dividend, // @[:@21494.4]
  input  [31:0] io_divisor, // @[:@21494.4]
  output [31:0] io_out // @[:@21494.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@21496.4]
  wire [29:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@21512.4]
  div_32_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@21496.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[31:2]; // @[ZynqBlackBoxes.scala 34:37:@21512.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@21513.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@21510.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@21509.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@21508.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@21507.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@21506.4 ZynqBlackBoxes.scala 33:17:@21511.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@21505.4]
endmodule
module x242_div( // @[:@21551.2]
  input         clock, // @[:@21552.4]
  input  [31:0] io_a, // @[:@21554.4]
  input         io_flow, // @[:@21554.4]
  output [31:0] io_result // @[:@21554.4]
);
  wire  x242_div_clock; // @[BigIPZynq.scala 25:21:@21562.4]
  wire  x242_div_io_flow; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] x242_div_io_dividend; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] x242_div_io_divisor; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] x242_div_io_out; // @[BigIPZynq.scala 25:21:@21562.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@21575.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@21575.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@21560.4]
  wire [31:0] _T_19; // @[BigIPZynq.scala 29:16:@21570.4]
  Divider x242_div ( // @[BigIPZynq.scala 25:21:@21562.4]
    .clock(x242_div_clock),
    .io_flow(x242_div_io_flow),
    .io_dividend(x242_div_io_dividend),
    .io_divisor(x242_div_io_divisor),
    .io_out(x242_div_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@21575.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@21560.4]
  assign _T_19 = $signed(x242_div_io_out); // @[BigIPZynq.scala 29:16:@21570.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@21583.4]
  assign x242_div_clock = clock; // @[:@21563.4]
  assign x242_div_io_flow = io_flow; // @[BigIPZynq.scala 28:17:@21569.4]
  assign x242_div_io_dividend = $unsigned(_T_15); // @[BigIPZynq.scala 26:21:@21566.4]
  assign x242_div_io_divisor = 32'h3; // @[BigIPZynq.scala 27:20:@21568.4]
  assign __io_b = $unsigned(_T_19); // @[Math.scala 721:17:@21578.4]
endmodule
module RetimeWrapper_243( // @[:@21597.2]
  input         clock, // @[:@21598.4]
  input         reset, // @[:@21599.4]
  input         io_flow, // @[:@21600.4]
  input  [31:0] io_in, // @[:@21600.4]
  output [31:0] io_out // @[:@21600.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21602.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@21602.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21615.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21614.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21613.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21612.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21611.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21609.4]
endmodule
module RetimeWrapper_245( // @[:@21808.2]
  input         clock, // @[:@21809.4]
  input         reset, // @[:@21810.4]
  input         io_flow, // @[:@21811.4]
  input  [31:0] io_in, // @[:@21811.4]
  output [31:0] io_out // @[:@21811.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21813.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@21813.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21826.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21825.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21824.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21823.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21822.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21820.4]
endmodule
module RetimeWrapper_246( // @[:@21840.2]
  input   clock, // @[:@21841.4]
  input   reset, // @[:@21842.4]
  input   io_flow, // @[:@21843.4]
  input   io_in, // @[:@21843.4]
  output  io_out // @[:@21843.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21845.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@21845.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21858.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21857.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@21856.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21855.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21854.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21852.4]
endmodule
module RetimeWrapper_247( // @[:@21872.2]
  input         clock, // @[:@21873.4]
  input         reset, // @[:@21874.4]
  input         io_flow, // @[:@21875.4]
  input  [31:0] io_in, // @[:@21875.4]
  output [31:0] io_out // @[:@21875.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21877.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21877.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21877.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21877.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21877.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21877.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@21877.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21890.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21889.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21888.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21887.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21886.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21884.4]
endmodule
module RetimeWrapper_249( // @[:@21936.2]
  input         clock, // @[:@21937.4]
  input         reset, // @[:@21938.4]
  input         io_flow, // @[:@21939.4]
  input  [31:0] io_in, // @[:@21939.4]
  output [31:0] io_out // @[:@21939.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21941.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@21941.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21954.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21953.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21952.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21951.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21950.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21948.4]
endmodule
module RetimeWrapper_251( // @[:@22000.2]
  input         clock, // @[:@22001.4]
  input         reset, // @[:@22002.4]
  input         io_flow, // @[:@22003.4]
  input  [31:0] io_in, // @[:@22003.4]
  output [31:0] io_out // @[:@22003.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22005.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@22005.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22018.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22017.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22016.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22015.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22014.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22012.4]
endmodule
module RetimeWrapper_256( // @[:@22160.2]
  input         clock, // @[:@22161.4]
  input         reset, // @[:@22162.4]
  input         io_flow, // @[:@22163.4]
  input  [31:0] io_in, // @[:@22163.4]
  output [31:0] io_out // @[:@22163.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22165.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@22165.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22178.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22177.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22176.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22175.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22174.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22172.4]
endmodule
module RetimeWrapper_257( // @[:@22192.2]
  input         clock, // @[:@22193.4]
  input         reset, // @[:@22194.4]
  input         io_flow, // @[:@22195.4]
  input  [31:0] io_in, // @[:@22195.4]
  output [31:0] io_out // @[:@22195.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22197.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@22197.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22210.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22209.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22208.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22207.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22206.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22204.4]
endmodule
module RetimeWrapper_258( // @[:@22224.2]
  input   clock, // @[:@22225.4]
  input   reset, // @[:@22226.4]
  input   io_flow, // @[:@22227.4]
  input   io_in, // @[:@22227.4]
  output  io_out // @[:@22227.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@22229.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@22229.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@22229.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22229.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22229.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22229.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@22229.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22242.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22241.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@22240.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22239.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22238.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22236.4]
endmodule
module RetimeWrapper_260( // @[:@22288.2]
  input         clock, // @[:@22289.4]
  input         reset, // @[:@22290.4]
  input         io_flow, // @[:@22291.4]
  input  [31:0] io_in, // @[:@22291.4]
  output [31:0] io_out // @[:@22291.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22293.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(37)) sr ( // @[RetimeShiftRegister.scala 15:20:@22293.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22306.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22305.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22304.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22303.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22302.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22300.4]
endmodule
module RetimeWrapper_277( // @[:@24117.2]
  input         clock, // @[:@24118.4]
  input         reset, // @[:@24119.4]
  input         io_flow, // @[:@24120.4]
  input  [31:0] io_in, // @[:@24120.4]
  output [31:0] io_out // @[:@24120.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24122.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(43)) sr ( // @[RetimeShiftRegister.scala 15:20:@24122.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24135.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24134.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@24133.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24132.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24131.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24129.4]
endmodule
module RetimeWrapper_279( // @[:@24328.2]
  input   clock, // @[:@24329.4]
  input   reset, // @[:@24330.4]
  input   io_flow, // @[:@24331.4]
  input   io_in, // @[:@24331.4]
  output  io_out // @[:@24331.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@24333.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@24333.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@24333.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24333.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24333.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24333.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@24333.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24346.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24345.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@24344.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24343.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24342.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24340.4]
endmodule
module RetimeWrapper_307( // @[:@26951.2]
  input         clock, // @[:@26952.4]
  input         reset, // @[:@26953.4]
  input         io_flow, // @[:@26954.4]
  input  [31:0] io_in, // @[:@26954.4]
  output [31:0] io_out // @[:@26954.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26956.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@26956.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26969.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26968.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26967.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26966.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26965.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26963.4]
endmodule
module RetimeWrapper_313( // @[:@27290.2]
  input         clock, // @[:@27291.4]
  input         reset, // @[:@27292.4]
  input         io_flow, // @[:@27293.4]
  input  [31:0] io_in, // @[:@27293.4]
  output [31:0] io_out // @[:@27293.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27295.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@27295.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27308.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27307.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27306.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27305.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27304.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27302.4]
endmodule
module Multiplier( // @[:@29118.2]
  input         clock, // @[:@29119.4]
  input         io_flow, // @[:@29121.4]
  input  [31:0] io_a, // @[:@29121.4]
  input  [31:0] io_b, // @[:@29121.4]
  output [31:0] io_out // @[:@29121.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@29123.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@29123.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@29123.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@29123.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@29123.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@29123.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@29133.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@29131.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@29130.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@29132.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@29129.4]
endmodule
module x312( // @[:@29153.2]
  input         clock, // @[:@29154.4]
  input  [31:0] io_a, // @[:@29156.4]
  input  [31:0] io_b, // @[:@29156.4]
  input         io_flow, // @[:@29156.4]
  output [31:0] io_result // @[:@29156.4]
);
  wire  x312_clock; // @[BigIPZynq.scala 63:21:@29163.4]
  wire  x312_io_flow; // @[BigIPZynq.scala 63:21:@29163.4]
  wire [31:0] x312_io_a; // @[BigIPZynq.scala 63:21:@29163.4]
  wire [31:0] x312_io_b; // @[BigIPZynq.scala 63:21:@29163.4]
  wire [31:0] x312_io_out; // @[BigIPZynq.scala 63:21:@29163.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@29172.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@29172.4]
  Multiplier x312 ( // @[BigIPZynq.scala 63:21:@29163.4]
    .clock(x312_clock),
    .io_flow(x312_io_flow),
    .io_a(x312_io_a),
    .io_b(x312_io_b),
    .io_out(x312_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@29172.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@29180.4]
  assign x312_clock = clock; // @[:@29164.4]
  assign x312_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@29168.4]
  assign x312_io_a = io_a; // @[BigIPZynq.scala 64:14:@29166.4]
  assign x312_io_b = io_b; // @[BigIPZynq.scala 65:14:@29167.4]
  assign fix2fixBox_io_a = x312_io_out; // @[Math.scala 254:23:@29175.4]
endmodule
module fix2fixBox_137( // @[:@29774.2]
  input  [31:0] io_a, // @[:@29777.4]
  output [32:0] io_b // @[:@29777.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@29791.4]
endmodule
module __87( // @[:@29793.2]
  input  [31:0] io_b, // @[:@29796.4]
  output [32:0] io_result // @[:@29796.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@29801.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@29801.4]
  fix2fixBox_137 fix2fixBox ( // @[BigIPZynq.scala 219:30:@29801.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@29809.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@29804.4]
endmodule
module x321_x7( // @[:@29905.2]
  input         clock, // @[:@29906.4]
  input         reset, // @[:@29907.4]
  input  [31:0] io_a, // @[:@29908.4]
  input  [31:0] io_b, // @[:@29908.4]
  input         io_flow, // @[:@29908.4]
  output [31:0] io_result // @[:@29908.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@29916.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@29916.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@29923.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@29923.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@29933.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@29933.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@29933.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@29933.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@29933.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@29921.4 Math.scala 724:14:@29922.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@29928.4 Math.scala 724:14:@29929.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@29930.4]
  __87 _ ( // @[Math.scala 720:24:@29916.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __87 __1 ( // @[Math.scala 720:24:@29923.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@29933.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@29921.4 Math.scala 724:14:@29922.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@29928.4 Math.scala 724:14:@29929.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@29930.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@29941.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@29919.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@29926.4]
  assign fix2fixBox_clock = clock; // @[:@29934.4]
  assign fix2fixBox_reset = reset; // @[:@29935.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@29936.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@29939.4]
endmodule
module RetimeWrapper_345( // @[:@30969.2]
  input         clock, // @[:@30970.4]
  input         reset, // @[:@30971.4]
  input         io_flow, // @[:@30972.4]
  input  [31:0] io_in, // @[:@30972.4]
  output [31:0] io_out // @[:@30972.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30974.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30974.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30974.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30974.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30974.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30974.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@30974.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30987.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30986.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30985.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30984.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30983.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30981.4]
endmodule
module fix2fixBox_161( // @[:@31158.2]
  input  [31:0] io_a, // @[:@31161.4]
  output [31:0] io_b // @[:@31161.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@31171.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@31171.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@31174.4]
endmodule
module x329( // @[:@31176.2]
  input  [31:0] io_b, // @[:@31179.4]
  output [31:0] io_result // @[:@31179.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@31184.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@31184.4]
  fix2fixBox_161 fix2fixBox ( // @[BigIPZynq.scala 219:30:@31184.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@31192.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@31187.4]
endmodule
module Multiplier_9( // @[:@31204.2]
  input         clock, // @[:@31205.4]
  input         io_flow, // @[:@31207.4]
  input  [38:0] io_a, // @[:@31207.4]
  input  [38:0] io_b, // @[:@31207.4]
  output [38:0] io_out // @[:@31207.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@31209.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@31209.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@31209.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@31209.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@31209.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@31209.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@31219.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@31217.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@31216.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@31218.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@31215.4]
endmodule
module fix2fixBox_162( // @[:@31221.2]
  input  [38:0] io_a, // @[:@31224.4]
  output [31:0] io_b // @[:@31224.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@31232.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@31235.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@31232.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@31235.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@31238.4]
endmodule
module x330_mul( // @[:@31240.2]
  input         clock, // @[:@31241.4]
  input  [31:0] io_a, // @[:@31243.4]
  input  [31:0] io_b, // @[:@31243.4]
  input         io_flow, // @[:@31243.4]
  output [31:0] io_result // @[:@31243.4]
);
  wire  x330_mul_clock; // @[BigIPZynq.scala 63:21:@31258.4]
  wire  x330_mul_io_flow; // @[BigIPZynq.scala 63:21:@31258.4]
  wire [38:0] x330_mul_io_a; // @[BigIPZynq.scala 63:21:@31258.4]
  wire [38:0] x330_mul_io_b; // @[BigIPZynq.scala 63:21:@31258.4]
  wire [38:0] x330_mul_io_out; // @[BigIPZynq.scala 63:21:@31258.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@31266.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@31266.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@31250.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@31252.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@31254.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@31256.4]
  Multiplier_9 x330_mul ( // @[BigIPZynq.scala 63:21:@31258.4]
    .clock(x330_mul_clock),
    .io_flow(x330_mul_io_flow),
    .io_a(x330_mul_io_a),
    .io_b(x330_mul_io_b),
    .io_out(x330_mul_io_out)
  );
  fix2fixBox_162 fix2fixBox ( // @[Math.scala 253:30:@31266.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@31250.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@31252.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@31254.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@31256.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@31274.4]
  assign x330_mul_clock = clock; // @[:@31259.4]
  assign x330_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@31263.4]
  assign x330_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@31261.4]
  assign x330_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@31262.4]
  assign fix2fixBox_io_a = x330_mul_io_out; // @[Math.scala 254:23:@31269.4]
endmodule
module fix2fixBox_163( // @[:@31276.2]
  input  [31:0] io_a, // @[:@31279.4]
  output [31:0] io_b // @[:@31279.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@31291.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@31291.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@31294.4]
endmodule
module x331( // @[:@31296.2]
  input  [31:0] io_b, // @[:@31299.4]
  output [31:0] io_result // @[:@31299.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@31304.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@31304.4]
  fix2fixBox_163 fix2fixBox ( // @[BigIPZynq.scala 219:30:@31304.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@31312.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@31307.4]
endmodule
module RetimeWrapper_347( // @[:@31326.2]
  input         clock, // @[:@31327.4]
  input         reset, // @[:@31328.4]
  input         io_flow, // @[:@31329.4]
  input  [31:0] io_in, // @[:@31329.4]
  output [31:0] io_out // @[:@31329.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31331.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31331.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31331.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31331.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31331.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31331.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(64)) sr ( // @[RetimeShiftRegister.scala 15:20:@31331.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31344.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31343.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31342.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31341.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31340.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31338.4]
endmodule
module RetimeWrapper_349( // @[:@31390.2]
  input   clock, // @[:@31391.4]
  input   reset, // @[:@31392.4]
  input   io_flow, // @[:@31393.4]
  input   io_in, // @[:@31393.4]
  output  io_out // @[:@31393.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@31395.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@31395.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@31395.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31395.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31395.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31395.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(64)) sr ( // @[RetimeShiftRegister.scala 15:20:@31395.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31408.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31407.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@31406.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31405.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31404.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31402.4]
endmodule
module RetimeWrapper_352( // @[:@31486.2]
  input         clock, // @[:@31487.4]
  input         reset, // @[:@31488.4]
  input         io_flow, // @[:@31489.4]
  input  [31:0] io_in, // @[:@31489.4]
  output [31:0] io_out // @[:@31489.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31491.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31491.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31491.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31491.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31491.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31491.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(56)) sr ( // @[RetimeShiftRegister.scala 15:20:@31491.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31504.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31503.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31502.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31501.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31500.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31498.4]
endmodule
module RetimeWrapper_354( // @[:@31550.2]
  input   clock, // @[:@31551.4]
  input   reset, // @[:@31552.4]
  input   io_flow, // @[:@31553.4]
  input   io_in, // @[:@31553.4]
  output  io_out // @[:@31553.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@31555.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@31555.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@31555.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31555.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31555.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31555.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(41)) sr ( // @[RetimeShiftRegister.scala 15:20:@31555.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31568.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31567.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@31566.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31565.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31564.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31562.4]
endmodule
module RetimeWrapper_355( // @[:@31582.2]
  input         clock, // @[:@31583.4]
  input         reset, // @[:@31584.4]
  input         io_flow, // @[:@31585.4]
  input  [31:0] io_in, // @[:@31585.4]
  output [31:0] io_out // @[:@31585.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31587.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31587.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31587.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31587.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31587.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31587.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(65)) sr ( // @[RetimeShiftRegister.scala 15:20:@31587.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31600.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31599.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31598.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31597.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31596.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31594.4]
endmodule
module RetimeWrapper_356( // @[:@31614.2]
  input         clock, // @[:@31615.4]
  input         reset, // @[:@31616.4]
  input         io_flow, // @[:@31617.4]
  input  [31:0] io_in, // @[:@31617.4]
  output [31:0] io_out // @[:@31617.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31619.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31619.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31619.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31619.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31619.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31619.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(44)) sr ( // @[RetimeShiftRegister.scala 15:20:@31619.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31632.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31631.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31630.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31629.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31628.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31626.4]
endmodule
module RetimeWrapper_357( // @[:@31646.2]
  input   clock, // @[:@31647.4]
  input   reset, // @[:@31648.4]
  input   io_flow, // @[:@31649.4]
  input   io_in, // @[:@31649.4]
  output  io_out // @[:@31649.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@31651.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@31651.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@31651.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31651.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31651.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31651.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(65)) sr ( // @[RetimeShiftRegister.scala 15:20:@31651.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31664.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31663.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@31662.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31661.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31660.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31658.4]
endmodule
module RetimeWrapper_359( // @[:@31710.2]
  input         clock, // @[:@31711.4]
  input         reset, // @[:@31712.4]
  input         io_flow, // @[:@31713.4]
  input  [31:0] io_in, // @[:@31713.4]
  output [31:0] io_out // @[:@31713.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31715.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31715.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31715.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31715.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31715.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31715.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(57)) sr ( // @[RetimeShiftRegister.scala 15:20:@31715.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31728.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31727.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31726.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31725.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31724.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31722.4]
endmodule
module RetimeWrapper_361( // @[:@31774.2]
  input   clock, // @[:@31775.4]
  input   reset, // @[:@31776.4]
  input   io_flow, // @[:@31777.4]
  input   io_in, // @[:@31777.4]
  output  io_out // @[:@31777.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@31779.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@31779.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@31779.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31779.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31779.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31779.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@31779.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31792.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31791.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@31790.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31789.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31788.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31786.4]
endmodule
module RetimeWrapper_362( // @[:@31806.2]
  input         clock, // @[:@31807.4]
  input         reset, // @[:@31808.4]
  input         io_flow, // @[:@31809.4]
  input  [31:0] io_in, // @[:@31809.4]
  output [31:0] io_out // @[:@31809.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31811.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31811.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31811.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31811.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31811.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31811.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(33)) sr ( // @[RetimeShiftRegister.scala 15:20:@31811.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31824.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31823.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31822.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31821.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31820.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31818.4]
endmodule
module RetimeWrapper_367( // @[:@31966.2]
  input         clock, // @[:@31967.4]
  input         reset, // @[:@31968.4]
  input         io_flow, // @[:@31969.4]
  input  [31:0] io_in, // @[:@31969.4]
  output [31:0] io_out // @[:@31969.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31971.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31971.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31971.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31971.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31971.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31971.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@31971.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31984.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31983.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31982.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31981.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31980.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31978.4]
endmodule
module RetimeWrapper_376( // @[:@33117.2]
  input   clock, // @[:@33118.4]
  input   reset, // @[:@33119.4]
  input   io_flow, // @[:@33120.4]
  input   io_in, // @[:@33120.4]
  output  io_out // @[:@33120.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@33122.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@33122.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@33122.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@33122.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@33122.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@33122.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(84)) sr ( // @[RetimeShiftRegister.scala 15:20:@33122.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@33135.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@33134.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@33133.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@33132.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@33131.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@33129.4]
endmodule
module x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@33201.2]
  input          clock, // @[:@33202.4]
  input          reset, // @[:@33203.4]
  output         io_in_x202_TVALID, // @[:@33204.4]
  input          io_in_x202_TREADY, // @[:@33204.4]
  output [255:0] io_in_x202_TDATA, // @[:@33204.4]
  output         io_in_x201_TREADY, // @[:@33204.4]
  input  [255:0] io_in_x201_TDATA, // @[:@33204.4]
  input  [7:0]   io_in_x201_TID, // @[:@33204.4]
  input  [7:0]   io_in_x201_TDEST, // @[:@33204.4]
  input          io_sigsIn_backpressure, // @[:@33204.4]
  input          io_sigsIn_datapathEn, // @[:@33204.4]
  input          io_sigsIn_break, // @[:@33204.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@33204.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@33204.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@33204.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@33204.4]
  input          io_rr // @[:@33204.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@33218.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@33218.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@33230.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@33230.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33253.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33253.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33253.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@33253.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@33253.4]
  wire  x233_lb_0_clock; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_reset; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_8_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_8_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_8_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_8_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_8_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_8_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_7_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_7_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_7_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_7_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_7_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_7_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_6_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_6_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_6_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_6_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_6_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_6_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_5_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_5_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_5_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_5_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_5_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_5_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_4_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_4_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_4_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_4_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_4_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_4_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_3_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_3_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_3_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_3_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_3_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_3_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_2_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_2_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_2_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_2_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_2_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_2_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_1_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_1_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_1_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_1_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_1_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_1_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_rPort_0_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_rPort_0_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_rPort_0_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_0_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_rPort_0_backpressure; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_rPort_0_output_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [1:0] x233_lb_0_io_wPort_0_banks_1; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [2:0] x233_lb_0_io_wPort_0_banks_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [9:0] x233_lb_0_io_wPort_0_ofs_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire [31:0] x233_lb_0_io_wPort_0_data_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x233_lb_0_io_wPort_0_en_0; // @[m_x233_lb_0.scala 35:17:@33263.4]
  wire  x234_lb2_0_clock; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_reset; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [1:0] x234_lb2_0_io_rPort_3_banks_1; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [2:0] x234_lb2_0_io_rPort_3_banks_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [9:0] x234_lb2_0_io_rPort_3_ofs_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_3_en_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_3_backpressure; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [31:0] x234_lb2_0_io_rPort_3_output_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [1:0] x234_lb2_0_io_rPort_2_banks_1; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [2:0] x234_lb2_0_io_rPort_2_banks_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [9:0] x234_lb2_0_io_rPort_2_ofs_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_2_en_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_2_backpressure; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [31:0] x234_lb2_0_io_rPort_2_output_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [1:0] x234_lb2_0_io_rPort_1_banks_1; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [2:0] x234_lb2_0_io_rPort_1_banks_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [9:0] x234_lb2_0_io_rPort_1_ofs_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_1_en_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_1_backpressure; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [31:0] x234_lb2_0_io_rPort_1_output_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [1:0] x234_lb2_0_io_rPort_0_banks_1; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [2:0] x234_lb2_0_io_rPort_0_banks_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [9:0] x234_lb2_0_io_rPort_0_ofs_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_0_en_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_rPort_0_backpressure; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [31:0] x234_lb2_0_io_rPort_0_output_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [1:0] x234_lb2_0_io_wPort_0_banks_1; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [2:0] x234_lb2_0_io_wPort_0_banks_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [9:0] x234_lb2_0_io_wPort_0_ofs_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire [31:0] x234_lb2_0_io_wPort_0_data_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x234_lb2_0_io_wPort_0_en_0; // @[m_x234_lb2_0.scala 30:17:@33330.4]
  wire  x414_sum_1_clock; // @[Math.scala 150:24:@33425.4]
  wire  x414_sum_1_reset; // @[Math.scala 150:24:@33425.4]
  wire [31:0] x414_sum_1_io_a; // @[Math.scala 150:24:@33425.4]
  wire [31:0] x414_sum_1_io_b; // @[Math.scala 150:24:@33425.4]
  wire  x414_sum_1_io_flow; // @[Math.scala 150:24:@33425.4]
  wire [31:0] x414_sum_1_io_result; // @[Math.scala 150:24:@33425.4]
  wire  x417_sum_1_clock; // @[Math.scala 150:24:@33463.4]
  wire  x417_sum_1_reset; // @[Math.scala 150:24:@33463.4]
  wire [31:0] x417_sum_1_io_a; // @[Math.scala 150:24:@33463.4]
  wire [31:0] x417_sum_1_io_b; // @[Math.scala 150:24:@33463.4]
  wire  x417_sum_1_io_flow; // @[Math.scala 150:24:@33463.4]
  wire [31:0] x417_sum_1_io_result; // @[Math.scala 150:24:@33463.4]
  wire  x420_sum_1_clock; // @[Math.scala 150:24:@33501.4]
  wire  x420_sum_1_reset; // @[Math.scala 150:24:@33501.4]
  wire [31:0] x420_sum_1_io_a; // @[Math.scala 150:24:@33501.4]
  wire [31:0] x420_sum_1_io_b; // @[Math.scala 150:24:@33501.4]
  wire  x420_sum_1_io_flow; // @[Math.scala 150:24:@33501.4]
  wire [31:0] x420_sum_1_io_result; // @[Math.scala 150:24:@33501.4]
  wire  x423_sum_1_clock; // @[Math.scala 150:24:@33539.4]
  wire  x423_sum_1_reset; // @[Math.scala 150:24:@33539.4]
  wire [31:0] x423_sum_1_io_a; // @[Math.scala 150:24:@33539.4]
  wire [31:0] x423_sum_1_io_b; // @[Math.scala 150:24:@33539.4]
  wire  x423_sum_1_io_flow; // @[Math.scala 150:24:@33539.4]
  wire [31:0] x423_sum_1_io_result; // @[Math.scala 150:24:@33539.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33562.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33562.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33562.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@33562.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@33562.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@33580.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@33580.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@33580.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@33580.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@33580.4]
  wire  x426_sum_1_clock; // @[Math.scala 150:24:@33593.4]
  wire  x426_sum_1_reset; // @[Math.scala 150:24:@33593.4]
  wire [31:0] x426_sum_1_io_a; // @[Math.scala 150:24:@33593.4]
  wire [31:0] x426_sum_1_io_b; // @[Math.scala 150:24:@33593.4]
  wire  x426_sum_1_io_flow; // @[Math.scala 150:24:@33593.4]
  wire [31:0] x426_sum_1_io_result; // @[Math.scala 150:24:@33593.4]
  wire  x429_sum_1_clock; // @[Math.scala 150:24:@33631.4]
  wire  x429_sum_1_reset; // @[Math.scala 150:24:@33631.4]
  wire [31:0] x429_sum_1_io_a; // @[Math.scala 150:24:@33631.4]
  wire [31:0] x429_sum_1_io_b; // @[Math.scala 150:24:@33631.4]
  wire  x429_sum_1_io_flow; // @[Math.scala 150:24:@33631.4]
  wire [31:0] x429_sum_1_io_result; // @[Math.scala 150:24:@33631.4]
  wire  x432_sub_1_clock; // @[Math.scala 191:24:@33657.4]
  wire  x432_sub_1_reset; // @[Math.scala 191:24:@33657.4]
  wire [31:0] x432_sub_1_io_a; // @[Math.scala 191:24:@33657.4]
  wire [31:0] x432_sub_1_io_b; // @[Math.scala 191:24:@33657.4]
  wire  x432_sub_1_io_flow; // @[Math.scala 191:24:@33657.4]
  wire [31:0] x432_sub_1_io_result; // @[Math.scala 191:24:@33657.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@33667.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@33667.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@33667.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@33667.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@33667.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@33676.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@33676.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@33676.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@33676.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@33676.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@33685.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@33685.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@33685.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@33685.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@33685.4]
  wire  x436_sum_1_clock; // @[Math.scala 150:24:@33724.4]
  wire  x436_sum_1_reset; // @[Math.scala 150:24:@33724.4]
  wire [31:0] x436_sum_1_io_a; // @[Math.scala 150:24:@33724.4]
  wire [31:0] x436_sum_1_io_b; // @[Math.scala 150:24:@33724.4]
  wire  x436_sum_1_io_flow; // @[Math.scala 150:24:@33724.4]
  wire [31:0] x436_sum_1_io_result; // @[Math.scala 150:24:@33724.4]
  wire  x242_div_1_clock; // @[Math.scala 327:24:@33736.4]
  wire [31:0] x242_div_1_io_a; // @[Math.scala 327:24:@33736.4]
  wire  x242_div_1_io_flow; // @[Math.scala 327:24:@33736.4]
  wire [31:0] x242_div_1_io_result; // @[Math.scala 327:24:@33736.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@33746.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@33746.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@33746.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@33746.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@33746.4]
  wire  x243_sum_1_clock; // @[Math.scala 150:24:@33755.4]
  wire  x243_sum_1_reset; // @[Math.scala 150:24:@33755.4]
  wire [31:0] x243_sum_1_io_a; // @[Math.scala 150:24:@33755.4]
  wire [31:0] x243_sum_1_io_b; // @[Math.scala 150:24:@33755.4]
  wire  x243_sum_1_io_flow; // @[Math.scala 150:24:@33755.4]
  wire [31:0] x243_sum_1_io_result; // @[Math.scala 150:24:@33755.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@33765.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@33765.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@33765.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@33774.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@33774.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@33774.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@33774.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@33774.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@33783.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@33783.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@33783.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@33783.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@33783.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@33792.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@33792.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@33792.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@33792.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@33792.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@33801.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@33801.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@33801.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@33801.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@33801.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@33833.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@33833.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@33833.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@33833.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@33833.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@33849.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@33849.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@33849.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@33849.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@33849.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@33858.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@33858.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@33858.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@33858.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@33858.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@33872.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@33872.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@33872.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@33872.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@33872.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@33887.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@33887.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@33887.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@33887.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@33887.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@33896.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@33896.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@33896.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@33896.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@33896.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@33905.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@33905.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@33905.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@33905.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@33905.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@33932.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@33932.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@33944.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@33944.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@33944.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@33944.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@33944.4]
  wire  x252_rdcol_1_clock; // @[Math.scala 191:24:@33967.4]
  wire  x252_rdcol_1_reset; // @[Math.scala 191:24:@33967.4]
  wire [31:0] x252_rdcol_1_io_a; // @[Math.scala 191:24:@33967.4]
  wire [31:0] x252_rdcol_1_io_b; // @[Math.scala 191:24:@33967.4]
  wire  x252_rdcol_1_io_flow; // @[Math.scala 191:24:@33967.4]
  wire [31:0] x252_rdcol_1_io_result; // @[Math.scala 191:24:@33967.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@33982.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@33982.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@33982.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@33982.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@33982.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@33991.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@33991.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@33991.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@33991.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@33991.4]
  wire  x439_sum_1_clock; // @[Math.scala 150:24:@34034.4]
  wire  x439_sum_1_reset; // @[Math.scala 150:24:@34034.4]
  wire [31:0] x439_sum_1_io_a; // @[Math.scala 150:24:@34034.4]
  wire [31:0] x439_sum_1_io_b; // @[Math.scala 150:24:@34034.4]
  wire  x439_sum_1_io_flow; // @[Math.scala 150:24:@34034.4]
  wire [31:0] x439_sum_1_io_result; // @[Math.scala 150:24:@34034.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@34057.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@34057.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@34057.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@34057.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@34057.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@34075.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@34075.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@34075.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@34075.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@34075.4]
  wire  x442_sum_1_clock; // @[Math.scala 150:24:@34088.4]
  wire  x442_sum_1_reset; // @[Math.scala 150:24:@34088.4]
  wire [31:0] x442_sum_1_io_a; // @[Math.scala 150:24:@34088.4]
  wire [31:0] x442_sum_1_io_b; // @[Math.scala 150:24:@34088.4]
  wire  x442_sum_1_io_flow; // @[Math.scala 150:24:@34088.4]
  wire [31:0] x442_sum_1_io_result; // @[Math.scala 150:24:@34088.4]
  wire  x445_sum_1_clock; // @[Math.scala 150:24:@34126.4]
  wire  x445_sum_1_reset; // @[Math.scala 150:24:@34126.4]
  wire [31:0] x445_sum_1_io_a; // @[Math.scala 150:24:@34126.4]
  wire [31:0] x445_sum_1_io_b; // @[Math.scala 150:24:@34126.4]
  wire  x445_sum_1_io_flow; // @[Math.scala 150:24:@34126.4]
  wire [31:0] x445_sum_1_io_result; // @[Math.scala 150:24:@34126.4]
  wire  x448_sum_1_clock; // @[Math.scala 150:24:@34164.4]
  wire  x448_sum_1_reset; // @[Math.scala 150:24:@34164.4]
  wire [31:0] x448_sum_1_io_a; // @[Math.scala 150:24:@34164.4]
  wire [31:0] x448_sum_1_io_b; // @[Math.scala 150:24:@34164.4]
  wire  x448_sum_1_io_flow; // @[Math.scala 150:24:@34164.4]
  wire [31:0] x448_sum_1_io_result; // @[Math.scala 150:24:@34164.4]
  wire  x451_sum_1_clock; // @[Math.scala 150:24:@34202.4]
  wire  x451_sum_1_reset; // @[Math.scala 150:24:@34202.4]
  wire [31:0] x451_sum_1_io_a; // @[Math.scala 150:24:@34202.4]
  wire [31:0] x451_sum_1_io_b; // @[Math.scala 150:24:@34202.4]
  wire  x451_sum_1_io_flow; // @[Math.scala 150:24:@34202.4]
  wire [31:0] x451_sum_1_io_result; // @[Math.scala 150:24:@34202.4]
  wire  x454_sum_1_clock; // @[Math.scala 150:24:@34240.4]
  wire  x454_sum_1_reset; // @[Math.scala 150:24:@34240.4]
  wire [31:0] x454_sum_1_io_a; // @[Math.scala 150:24:@34240.4]
  wire [31:0] x454_sum_1_io_b; // @[Math.scala 150:24:@34240.4]
  wire  x454_sum_1_io_flow; // @[Math.scala 150:24:@34240.4]
  wire [31:0] x454_sum_1_io_result; // @[Math.scala 150:24:@34240.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@34255.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@34255.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@34255.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@34255.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@34255.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@34269.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@34269.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@34269.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@34269.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@34269.4]
  wire  x457_sub_1_clock; // @[Math.scala 191:24:@34280.4]
  wire  x457_sub_1_reset; // @[Math.scala 191:24:@34280.4]
  wire [31:0] x457_sub_1_io_a; // @[Math.scala 191:24:@34280.4]
  wire [31:0] x457_sub_1_io_b; // @[Math.scala 191:24:@34280.4]
  wire  x457_sub_1_io_flow; // @[Math.scala 191:24:@34280.4]
  wire [31:0] x457_sub_1_io_result; // @[Math.scala 191:24:@34280.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@34290.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@34290.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@34290.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@34290.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@34290.4]
  wire  x257_div_1_clock; // @[Math.scala 327:24:@34304.4]
  wire [31:0] x257_div_1_io_a; // @[Math.scala 327:24:@34304.4]
  wire  x257_div_1_io_flow; // @[Math.scala 327:24:@34304.4]
  wire [31:0] x257_div_1_io_result; // @[Math.scala 327:24:@34304.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@34314.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@34314.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@34314.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@34314.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@34314.4]
  wire  x258_sum_1_clock; // @[Math.scala 150:24:@34323.4]
  wire  x258_sum_1_reset; // @[Math.scala 150:24:@34323.4]
  wire [31:0] x258_sum_1_io_a; // @[Math.scala 150:24:@34323.4]
  wire [31:0] x258_sum_1_io_b; // @[Math.scala 150:24:@34323.4]
  wire  x258_sum_1_io_flow; // @[Math.scala 150:24:@34323.4]
  wire [31:0] x258_sum_1_io_result; // @[Math.scala 150:24:@34323.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@34333.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@34333.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@34333.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@34333.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@34333.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@34342.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@34342.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@34342.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@34342.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@34342.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@34354.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@34354.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@34354.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@34354.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@34354.4]
  wire  x261_rdcol_1_clock; // @[Math.scala 191:24:@34377.4]
  wire  x261_rdcol_1_reset; // @[Math.scala 191:24:@34377.4]
  wire [31:0] x261_rdcol_1_io_a; // @[Math.scala 191:24:@34377.4]
  wire [31:0] x261_rdcol_1_io_b; // @[Math.scala 191:24:@34377.4]
  wire  x261_rdcol_1_io_flow; // @[Math.scala 191:24:@34377.4]
  wire [31:0] x261_rdcol_1_io_result; // @[Math.scala 191:24:@34377.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@34394.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@34394.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@34394.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@34394.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@34394.4]
  wire  x461_sum_1_clock; // @[Math.scala 150:24:@34437.4]
  wire  x461_sum_1_reset; // @[Math.scala 150:24:@34437.4]
  wire [31:0] x461_sum_1_io_a; // @[Math.scala 150:24:@34437.4]
  wire [31:0] x461_sum_1_io_b; // @[Math.scala 150:24:@34437.4]
  wire  x461_sum_1_io_flow; // @[Math.scala 150:24:@34437.4]
  wire [31:0] x461_sum_1_io_result; // @[Math.scala 150:24:@34437.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@34460.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@34460.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@34460.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@34460.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@34460.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@34478.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@34478.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@34478.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@34478.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@34478.4]
  wire  x464_sum_1_clock; // @[Math.scala 150:24:@34491.4]
  wire  x464_sum_1_reset; // @[Math.scala 150:24:@34491.4]
  wire [31:0] x464_sum_1_io_a; // @[Math.scala 150:24:@34491.4]
  wire [31:0] x464_sum_1_io_b; // @[Math.scala 150:24:@34491.4]
  wire  x464_sum_1_io_flow; // @[Math.scala 150:24:@34491.4]
  wire [31:0] x464_sum_1_io_result; // @[Math.scala 150:24:@34491.4]
  wire  x467_sum_1_clock; // @[Math.scala 150:24:@34529.4]
  wire  x467_sum_1_reset; // @[Math.scala 150:24:@34529.4]
  wire [31:0] x467_sum_1_io_a; // @[Math.scala 150:24:@34529.4]
  wire [31:0] x467_sum_1_io_b; // @[Math.scala 150:24:@34529.4]
  wire  x467_sum_1_io_flow; // @[Math.scala 150:24:@34529.4]
  wire [31:0] x467_sum_1_io_result; // @[Math.scala 150:24:@34529.4]
  wire  x470_sum_1_clock; // @[Math.scala 150:24:@34567.4]
  wire  x470_sum_1_reset; // @[Math.scala 150:24:@34567.4]
  wire [31:0] x470_sum_1_io_a; // @[Math.scala 150:24:@34567.4]
  wire [31:0] x470_sum_1_io_b; // @[Math.scala 150:24:@34567.4]
  wire  x470_sum_1_io_flow; // @[Math.scala 150:24:@34567.4]
  wire [31:0] x470_sum_1_io_result; // @[Math.scala 150:24:@34567.4]
  wire  x473_sum_1_clock; // @[Math.scala 150:24:@34605.4]
  wire  x473_sum_1_reset; // @[Math.scala 150:24:@34605.4]
  wire [31:0] x473_sum_1_io_a; // @[Math.scala 150:24:@34605.4]
  wire [31:0] x473_sum_1_io_b; // @[Math.scala 150:24:@34605.4]
  wire  x473_sum_1_io_flow; // @[Math.scala 150:24:@34605.4]
  wire [31:0] x473_sum_1_io_result; // @[Math.scala 150:24:@34605.4]
  wire  x476_sum_1_clock; // @[Math.scala 150:24:@34643.4]
  wire  x476_sum_1_reset; // @[Math.scala 150:24:@34643.4]
  wire [31:0] x476_sum_1_io_a; // @[Math.scala 150:24:@34643.4]
  wire [31:0] x476_sum_1_io_b; // @[Math.scala 150:24:@34643.4]
  wire  x476_sum_1_io_flow; // @[Math.scala 150:24:@34643.4]
  wire [31:0] x476_sum_1_io_result; // @[Math.scala 150:24:@34643.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@34658.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@34658.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@34658.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@34658.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@34658.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@34672.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@34672.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@34672.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@34672.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@34672.4]
  wire  x479_sub_1_clock; // @[Math.scala 191:24:@34683.4]
  wire  x479_sub_1_reset; // @[Math.scala 191:24:@34683.4]
  wire [31:0] x479_sub_1_io_a; // @[Math.scala 191:24:@34683.4]
  wire [31:0] x479_sub_1_io_b; // @[Math.scala 191:24:@34683.4]
  wire  x479_sub_1_io_flow; // @[Math.scala 191:24:@34683.4]
  wire [31:0] x479_sub_1_io_result; // @[Math.scala 191:24:@34683.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@34693.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@34693.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@34693.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@34693.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@34693.4]
  wire  x266_div_1_clock; // @[Math.scala 327:24:@34707.4]
  wire [31:0] x266_div_1_io_a; // @[Math.scala 327:24:@34707.4]
  wire  x266_div_1_io_flow; // @[Math.scala 327:24:@34707.4]
  wire [31:0] x266_div_1_io_result; // @[Math.scala 327:24:@34707.4]
  wire  x267_sum_1_clock; // @[Math.scala 150:24:@34717.4]
  wire  x267_sum_1_reset; // @[Math.scala 150:24:@34717.4]
  wire [31:0] x267_sum_1_io_a; // @[Math.scala 150:24:@34717.4]
  wire [31:0] x267_sum_1_io_b; // @[Math.scala 150:24:@34717.4]
  wire  x267_sum_1_io_flow; // @[Math.scala 150:24:@34717.4]
  wire [31:0] x267_sum_1_io_result; // @[Math.scala 150:24:@34717.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@34727.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@34727.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@34727.4]
  wire [31:0] RetimeWrapper_41_io_in; // @[package.scala 93:22:@34727.4]
  wire [31:0] RetimeWrapper_41_io_out; // @[package.scala 93:22:@34727.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@34736.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@34736.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@34736.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@34736.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@34736.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@34748.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@34748.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@34748.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@34748.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@34748.4]
  wire  x270_rdrow_1_clock; // @[Math.scala 191:24:@34771.4]
  wire  x270_rdrow_1_reset; // @[Math.scala 191:24:@34771.4]
  wire [31:0] x270_rdrow_1_io_a; // @[Math.scala 191:24:@34771.4]
  wire [31:0] x270_rdrow_1_io_b; // @[Math.scala 191:24:@34771.4]
  wire  x270_rdrow_1_io_flow; // @[Math.scala 191:24:@34771.4]
  wire [31:0] x270_rdrow_1_io_result; // @[Math.scala 191:24:@34771.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@34797.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@34797.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@34797.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@34797.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@34797.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@34806.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@34806.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@34806.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@34806.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@34806.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@34828.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@34828.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@34828.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@34828.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@34828.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@34854.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@34854.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@34854.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@34854.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@34854.4]
  wire  x485_sum_1_clock; // @[Math.scala 150:24:@34875.4]
  wire  x485_sum_1_reset; // @[Math.scala 150:24:@34875.4]
  wire [31:0] x485_sum_1_io_a; // @[Math.scala 150:24:@34875.4]
  wire [31:0] x485_sum_1_io_b; // @[Math.scala 150:24:@34875.4]
  wire  x485_sum_1_io_flow; // @[Math.scala 150:24:@34875.4]
  wire [31:0] x485_sum_1_io_result; // @[Math.scala 150:24:@34875.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@34885.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@34885.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@34885.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@34894.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@34894.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@34894.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@34894.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@34894.4]
  wire  x278_sum_1_clock; // @[Math.scala 150:24:@34903.4]
  wire  x278_sum_1_reset; // @[Math.scala 150:24:@34903.4]
  wire [31:0] x278_sum_1_io_a; // @[Math.scala 150:24:@34903.4]
  wire [31:0] x278_sum_1_io_b; // @[Math.scala 150:24:@34903.4]
  wire  x278_sum_1_io_flow; // @[Math.scala 150:24:@34903.4]
  wire [31:0] x278_sum_1_io_result; // @[Math.scala 150:24:@34903.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@34913.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@34913.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@34913.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@34913.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@34913.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@34922.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@34922.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@34931.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@34931.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@34931.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@34931.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@34931.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@34943.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@34943.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@34943.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@34943.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@34943.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@34970.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@34970.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@34970.4]
  wire  x283_sum_1_clock; // @[Math.scala 150:24:@34981.4]
  wire  x283_sum_1_reset; // @[Math.scala 150:24:@34981.4]
  wire [31:0] x283_sum_1_io_a; // @[Math.scala 150:24:@34981.4]
  wire [31:0] x283_sum_1_io_b; // @[Math.scala 150:24:@34981.4]
  wire  x283_sum_1_io_flow; // @[Math.scala 150:24:@34981.4]
  wire [31:0] x283_sum_1_io_result; // @[Math.scala 150:24:@34981.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@34991.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@34991.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@34991.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@34991.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@34991.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@35003.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@35003.4]
  wire  x288_sum_1_clock; // @[Math.scala 150:24:@35030.4]
  wire  x288_sum_1_reset; // @[Math.scala 150:24:@35030.4]
  wire [31:0] x288_sum_1_io_a; // @[Math.scala 150:24:@35030.4]
  wire [31:0] x288_sum_1_io_b; // @[Math.scala 150:24:@35030.4]
  wire  x288_sum_1_io_flow; // @[Math.scala 150:24:@35030.4]
  wire [31:0] x288_sum_1_io_result; // @[Math.scala 150:24:@35030.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@35052.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@35052.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@35052.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@35052.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@35052.4]
  wire  x291_rdrow_1_clock; // @[Math.scala 191:24:@35075.4]
  wire  x291_rdrow_1_reset; // @[Math.scala 191:24:@35075.4]
  wire [31:0] x291_rdrow_1_io_a; // @[Math.scala 191:24:@35075.4]
  wire [31:0] x291_rdrow_1_io_b; // @[Math.scala 191:24:@35075.4]
  wire  x291_rdrow_1_io_flow; // @[Math.scala 191:24:@35075.4]
  wire [31:0] x291_rdrow_1_io_result; // @[Math.scala 191:24:@35075.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@35101.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@35101.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@35101.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@35101.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@35101.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@35123.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@35123.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@35123.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@35123.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@35123.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@35149.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@35149.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@35149.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@35149.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@35149.4]
  wire  x490_sum_1_clock; // @[Math.scala 150:24:@35170.4]
  wire  x490_sum_1_reset; // @[Math.scala 150:24:@35170.4]
  wire [31:0] x490_sum_1_io_a; // @[Math.scala 150:24:@35170.4]
  wire [31:0] x490_sum_1_io_b; // @[Math.scala 150:24:@35170.4]
  wire  x490_sum_1_io_flow; // @[Math.scala 150:24:@35170.4]
  wire [31:0] x490_sum_1_io_result; // @[Math.scala 150:24:@35170.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@35180.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@35180.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@35180.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@35180.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@35180.4]
  wire  x299_sum_1_clock; // @[Math.scala 150:24:@35189.4]
  wire  x299_sum_1_reset; // @[Math.scala 150:24:@35189.4]
  wire [31:0] x299_sum_1_io_a; // @[Math.scala 150:24:@35189.4]
  wire [31:0] x299_sum_1_io_b; // @[Math.scala 150:24:@35189.4]
  wire  x299_sum_1_io_flow; // @[Math.scala 150:24:@35189.4]
  wire [31:0] x299_sum_1_io_result; // @[Math.scala 150:24:@35189.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@35199.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@35199.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@35199.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@35199.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@35199.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@35208.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@35208.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@35208.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@35208.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@35208.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@35217.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@35217.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@35217.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@35217.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@35217.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@35229.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@35229.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@35229.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@35229.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@35229.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@35256.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@35256.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@35256.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@35256.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@35256.4]
  wire  x304_sum_1_clock; // @[Math.scala 150:24:@35265.4]
  wire  x304_sum_1_reset; // @[Math.scala 150:24:@35265.4]
  wire [31:0] x304_sum_1_io_a; // @[Math.scala 150:24:@35265.4]
  wire [31:0] x304_sum_1_io_b; // @[Math.scala 150:24:@35265.4]
  wire  x304_sum_1_io_flow; // @[Math.scala 150:24:@35265.4]
  wire [31:0] x304_sum_1_io_result; // @[Math.scala 150:24:@35265.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@35275.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@35275.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@35275.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@35275.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@35275.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@35287.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@35287.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@35287.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@35287.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@35287.4]
  wire  x309_sum_1_clock; // @[Math.scala 150:24:@35314.4]
  wire  x309_sum_1_reset; // @[Math.scala 150:24:@35314.4]
  wire [31:0] x309_sum_1_io_a; // @[Math.scala 150:24:@35314.4]
  wire [31:0] x309_sum_1_io_b; // @[Math.scala 150:24:@35314.4]
  wire  x309_sum_1_io_flow; // @[Math.scala 150:24:@35314.4]
  wire [31:0] x309_sum_1_io_result; // @[Math.scala 150:24:@35314.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@35324.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@35324.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@35324.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@35324.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@35324.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@35336.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@35336.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@35336.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@35336.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@35336.4]
  wire  x312_1_clock; // @[Math.scala 262:24:@35359.4]
  wire [31:0] x312_1_io_a; // @[Math.scala 262:24:@35359.4]
  wire [31:0] x312_1_io_b; // @[Math.scala 262:24:@35359.4]
  wire  x312_1_io_flow; // @[Math.scala 262:24:@35359.4]
  wire [31:0] x312_1_io_result; // @[Math.scala 262:24:@35359.4]
  wire  x313_1_clock; // @[Math.scala 262:24:@35371.4]
  wire [31:0] x313_1_io_a; // @[Math.scala 262:24:@35371.4]
  wire [31:0] x313_1_io_b; // @[Math.scala 262:24:@35371.4]
  wire  x313_1_io_flow; // @[Math.scala 262:24:@35371.4]
  wire [31:0] x313_1_io_result; // @[Math.scala 262:24:@35371.4]
  wire  x314_1_clock; // @[Math.scala 262:24:@35383.4]
  wire [31:0] x314_1_io_a; // @[Math.scala 262:24:@35383.4]
  wire [31:0] x314_1_io_b; // @[Math.scala 262:24:@35383.4]
  wire  x314_1_io_flow; // @[Math.scala 262:24:@35383.4]
  wire [31:0] x314_1_io_result; // @[Math.scala 262:24:@35383.4]
  wire  x315_1_clock; // @[Math.scala 262:24:@35395.4]
  wire [31:0] x315_1_io_a; // @[Math.scala 262:24:@35395.4]
  wire [31:0] x315_1_io_b; // @[Math.scala 262:24:@35395.4]
  wire  x315_1_io_flow; // @[Math.scala 262:24:@35395.4]
  wire [31:0] x315_1_io_result; // @[Math.scala 262:24:@35395.4]
  wire  x316_1_clock; // @[Math.scala 262:24:@35409.4]
  wire [31:0] x316_1_io_a; // @[Math.scala 262:24:@35409.4]
  wire [31:0] x316_1_io_b; // @[Math.scala 262:24:@35409.4]
  wire  x316_1_io_flow; // @[Math.scala 262:24:@35409.4]
  wire [31:0] x316_1_io_result; // @[Math.scala 262:24:@35409.4]
  wire  x317_1_clock; // @[Math.scala 262:24:@35421.4]
  wire [31:0] x317_1_io_a; // @[Math.scala 262:24:@35421.4]
  wire [31:0] x317_1_io_b; // @[Math.scala 262:24:@35421.4]
  wire  x317_1_io_flow; // @[Math.scala 262:24:@35421.4]
  wire [31:0] x317_1_io_result; // @[Math.scala 262:24:@35421.4]
  wire  x318_1_clock; // @[Math.scala 262:24:@35433.4]
  wire [31:0] x318_1_io_a; // @[Math.scala 262:24:@35433.4]
  wire [31:0] x318_1_io_b; // @[Math.scala 262:24:@35433.4]
  wire  x318_1_io_flow; // @[Math.scala 262:24:@35433.4]
  wire [31:0] x318_1_io_result; // @[Math.scala 262:24:@35433.4]
  wire  x319_1_clock; // @[Math.scala 262:24:@35445.4]
  wire [31:0] x319_1_io_a; // @[Math.scala 262:24:@35445.4]
  wire [31:0] x319_1_io_b; // @[Math.scala 262:24:@35445.4]
  wire  x319_1_io_flow; // @[Math.scala 262:24:@35445.4]
  wire [31:0] x319_1_io_result; // @[Math.scala 262:24:@35445.4]
  wire  x320_1_clock; // @[Math.scala 262:24:@35457.4]
  wire [31:0] x320_1_io_a; // @[Math.scala 262:24:@35457.4]
  wire [31:0] x320_1_io_b; // @[Math.scala 262:24:@35457.4]
  wire  x320_1_io_flow; // @[Math.scala 262:24:@35457.4]
  wire [31:0] x320_1_io_result; // @[Math.scala 262:24:@35457.4]
  wire  x321_x7_1_clock; // @[Math.scala 150:24:@35467.4]
  wire  x321_x7_1_reset; // @[Math.scala 150:24:@35467.4]
  wire [31:0] x321_x7_1_io_a; // @[Math.scala 150:24:@35467.4]
  wire [31:0] x321_x7_1_io_b; // @[Math.scala 150:24:@35467.4]
  wire  x321_x7_1_io_flow; // @[Math.scala 150:24:@35467.4]
  wire [31:0] x321_x7_1_io_result; // @[Math.scala 150:24:@35467.4]
  wire  x322_x8_1_clock; // @[Math.scala 150:24:@35477.4]
  wire  x322_x8_1_reset; // @[Math.scala 150:24:@35477.4]
  wire [31:0] x322_x8_1_io_a; // @[Math.scala 150:24:@35477.4]
  wire [31:0] x322_x8_1_io_b; // @[Math.scala 150:24:@35477.4]
  wire  x322_x8_1_io_flow; // @[Math.scala 150:24:@35477.4]
  wire [31:0] x322_x8_1_io_result; // @[Math.scala 150:24:@35477.4]
  wire  x323_x7_1_clock; // @[Math.scala 150:24:@35487.4]
  wire  x323_x7_1_reset; // @[Math.scala 150:24:@35487.4]
  wire [31:0] x323_x7_1_io_a; // @[Math.scala 150:24:@35487.4]
  wire [31:0] x323_x7_1_io_b; // @[Math.scala 150:24:@35487.4]
  wire  x323_x7_1_io_flow; // @[Math.scala 150:24:@35487.4]
  wire [31:0] x323_x7_1_io_result; // @[Math.scala 150:24:@35487.4]
  wire  x324_x8_1_clock; // @[Math.scala 150:24:@35497.4]
  wire  x324_x8_1_reset; // @[Math.scala 150:24:@35497.4]
  wire [31:0] x324_x8_1_io_a; // @[Math.scala 150:24:@35497.4]
  wire [31:0] x324_x8_1_io_b; // @[Math.scala 150:24:@35497.4]
  wire  x324_x8_1_io_flow; // @[Math.scala 150:24:@35497.4]
  wire [31:0] x324_x8_1_io_result; // @[Math.scala 150:24:@35497.4]
  wire  x325_x7_1_clock; // @[Math.scala 150:24:@35507.4]
  wire  x325_x7_1_reset; // @[Math.scala 150:24:@35507.4]
  wire [31:0] x325_x7_1_io_a; // @[Math.scala 150:24:@35507.4]
  wire [31:0] x325_x7_1_io_b; // @[Math.scala 150:24:@35507.4]
  wire  x325_x7_1_io_flow; // @[Math.scala 150:24:@35507.4]
  wire [31:0] x325_x7_1_io_result; // @[Math.scala 150:24:@35507.4]
  wire  x326_x8_1_clock; // @[Math.scala 150:24:@35517.4]
  wire  x326_x8_1_reset; // @[Math.scala 150:24:@35517.4]
  wire [31:0] x326_x8_1_io_a; // @[Math.scala 150:24:@35517.4]
  wire [31:0] x326_x8_1_io_b; // @[Math.scala 150:24:@35517.4]
  wire  x326_x8_1_io_flow; // @[Math.scala 150:24:@35517.4]
  wire [31:0] x326_x8_1_io_result; // @[Math.scala 150:24:@35517.4]
  wire  x327_x7_1_clock; // @[Math.scala 150:24:@35527.4]
  wire  x327_x7_1_reset; // @[Math.scala 150:24:@35527.4]
  wire [31:0] x327_x7_1_io_a; // @[Math.scala 150:24:@35527.4]
  wire [31:0] x327_x7_1_io_b; // @[Math.scala 150:24:@35527.4]
  wire  x327_x7_1_io_flow; // @[Math.scala 150:24:@35527.4]
  wire [31:0] x327_x7_1_io_result; // @[Math.scala 150:24:@35527.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@35537.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@35537.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@35537.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@35537.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@35537.4]
  wire  x328_sum_1_clock; // @[Math.scala 150:24:@35546.4]
  wire  x328_sum_1_reset; // @[Math.scala 150:24:@35546.4]
  wire [31:0] x328_sum_1_io_a; // @[Math.scala 150:24:@35546.4]
  wire [31:0] x328_sum_1_io_b; // @[Math.scala 150:24:@35546.4]
  wire  x328_sum_1_io_flow; // @[Math.scala 150:24:@35546.4]
  wire [31:0] x328_sum_1_io_result; // @[Math.scala 150:24:@35546.4]
  wire [31:0] x329_1_io_b; // @[Math.scala 720:24:@35556.4]
  wire [31:0] x329_1_io_result; // @[Math.scala 720:24:@35556.4]
  wire  x330_mul_1_clock; // @[Math.scala 262:24:@35567.4]
  wire [31:0] x330_mul_1_io_a; // @[Math.scala 262:24:@35567.4]
  wire [31:0] x330_mul_1_io_b; // @[Math.scala 262:24:@35567.4]
  wire  x330_mul_1_io_flow; // @[Math.scala 262:24:@35567.4]
  wire [31:0] x330_mul_1_io_result; // @[Math.scala 262:24:@35567.4]
  wire [31:0] x331_1_io_b; // @[Math.scala 720:24:@35577.4]
  wire [31:0] x331_1_io_result; // @[Math.scala 720:24:@35577.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@35586.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@35586.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@35586.4]
  wire [31:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@35586.4]
  wire [31:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@35586.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@35595.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@35595.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@35595.4]
  wire [31:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@35595.4]
  wire [31:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@35595.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@35604.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@35604.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@35604.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@35604.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@35604.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@35613.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@35613.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@35613.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@35613.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@35613.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@35622.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@35622.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@35622.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@35622.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@35622.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@35631.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@35631.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@35631.4]
  wire [31:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@35631.4]
  wire [31:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@35631.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@35663.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@35663.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@35663.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@35663.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@35663.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@35672.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@35672.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@35672.4]
  wire [31:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@35672.4]
  wire [31:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@35672.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@35681.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@35681.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@35681.4]
  wire [31:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@35681.4]
  wire [31:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@35681.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@35699.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@35699.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@35699.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@35699.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@35699.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@35708.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@35708.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@35708.4]
  wire [31:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@35708.4]
  wire [31:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@35708.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@35720.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@35720.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@35720.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@35720.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@35720.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@35741.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@35741.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@35741.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@35741.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@35741.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@35750.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@35750.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@35750.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@35750.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@35750.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@35759.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@35759.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@35759.4]
  wire [31:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@35759.4]
  wire [31:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@35759.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@35771.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@35771.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@35771.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@35771.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@35771.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@35792.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@35792.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@35792.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@35792.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@35792.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@35801.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@35801.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@35801.4]
  wire [31:0] RetimeWrapper_92_io_in; // @[package.scala 93:22:@35801.4]
  wire [31:0] RetimeWrapper_92_io_out; // @[package.scala 93:22:@35801.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@35810.4]
  wire [31:0] RetimeWrapper_93_io_in; // @[package.scala 93:22:@35810.4]
  wire [31:0] RetimeWrapper_93_io_out; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@35822.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@35822.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@35822.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@35822.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@35822.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@35843.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@35843.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@35843.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@35843.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@35843.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@35852.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@35852.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@35852.4]
  wire [31:0] RetimeWrapper_96_io_in; // @[package.scala 93:22:@35852.4]
  wire [31:0] RetimeWrapper_96_io_out; // @[package.scala 93:22:@35852.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@35864.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@35864.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@35864.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@35864.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@35864.4]
  wire  x343_1_clock; // @[Math.scala 262:24:@35887.4]
  wire [31:0] x343_1_io_a; // @[Math.scala 262:24:@35887.4]
  wire [31:0] x343_1_io_b; // @[Math.scala 262:24:@35887.4]
  wire  x343_1_io_flow; // @[Math.scala 262:24:@35887.4]
  wire [31:0] x343_1_io_result; // @[Math.scala 262:24:@35887.4]
  wire  x344_1_clock; // @[Math.scala 262:24:@35901.4]
  wire [31:0] x344_1_io_a; // @[Math.scala 262:24:@35901.4]
  wire [31:0] x344_1_io_b; // @[Math.scala 262:24:@35901.4]
  wire  x344_1_io_flow; // @[Math.scala 262:24:@35901.4]
  wire [31:0] x344_1_io_result; // @[Math.scala 262:24:@35901.4]
  wire  x345_1_clock; // @[Math.scala 262:24:@35913.4]
  wire [31:0] x345_1_io_a; // @[Math.scala 262:24:@35913.4]
  wire [31:0] x345_1_io_b; // @[Math.scala 262:24:@35913.4]
  wire  x345_1_io_flow; // @[Math.scala 262:24:@35913.4]
  wire [31:0] x345_1_io_result; // @[Math.scala 262:24:@35913.4]
  wire  x346_1_clock; // @[Math.scala 262:24:@35925.4]
  wire [31:0] x346_1_io_a; // @[Math.scala 262:24:@35925.4]
  wire [31:0] x346_1_io_b; // @[Math.scala 262:24:@35925.4]
  wire  x346_1_io_flow; // @[Math.scala 262:24:@35925.4]
  wire [31:0] x346_1_io_result; // @[Math.scala 262:24:@35925.4]
  wire  x347_x9_1_clock; // @[Math.scala 150:24:@35935.4]
  wire  x347_x9_1_reset; // @[Math.scala 150:24:@35935.4]
  wire [31:0] x347_x9_1_io_a; // @[Math.scala 150:24:@35935.4]
  wire [31:0] x347_x9_1_io_b; // @[Math.scala 150:24:@35935.4]
  wire  x347_x9_1_io_flow; // @[Math.scala 150:24:@35935.4]
  wire [31:0] x347_x9_1_io_result; // @[Math.scala 150:24:@35935.4]
  wire  x348_x10_1_clock; // @[Math.scala 150:24:@35945.4]
  wire  x348_x10_1_reset; // @[Math.scala 150:24:@35945.4]
  wire [31:0] x348_x10_1_io_a; // @[Math.scala 150:24:@35945.4]
  wire [31:0] x348_x10_1_io_b; // @[Math.scala 150:24:@35945.4]
  wire  x348_x10_1_io_flow; // @[Math.scala 150:24:@35945.4]
  wire [31:0] x348_x10_1_io_result; // @[Math.scala 150:24:@35945.4]
  wire  x349_sum_1_clock; // @[Math.scala 150:24:@35955.4]
  wire  x349_sum_1_reset; // @[Math.scala 150:24:@35955.4]
  wire [31:0] x349_sum_1_io_a; // @[Math.scala 150:24:@35955.4]
  wire [31:0] x349_sum_1_io_b; // @[Math.scala 150:24:@35955.4]
  wire  x349_sum_1_io_flow; // @[Math.scala 150:24:@35955.4]
  wire [31:0] x349_sum_1_io_result; // @[Math.scala 150:24:@35955.4]
  wire [31:0] x350_1_io_b; // @[Math.scala 720:24:@35965.4]
  wire [31:0] x350_1_io_result; // @[Math.scala 720:24:@35965.4]
  wire  x351_mul_1_clock; // @[Math.scala 262:24:@35976.4]
  wire [31:0] x351_mul_1_io_a; // @[Math.scala 262:24:@35976.4]
  wire [31:0] x351_mul_1_io_b; // @[Math.scala 262:24:@35976.4]
  wire  x351_mul_1_io_flow; // @[Math.scala 262:24:@35976.4]
  wire [31:0] x351_mul_1_io_result; // @[Math.scala 262:24:@35976.4]
  wire [31:0] x352_1_io_b; // @[Math.scala 720:24:@35986.4]
  wire [31:0] x352_1_io_result; // @[Math.scala 720:24:@35986.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@35999.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@35999.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@35999.4]
  wire [31:0] RetimeWrapper_98_io_in; // @[package.scala 93:22:@35999.4]
  wire [31:0] RetimeWrapper_98_io_out; // @[package.scala 93:22:@35999.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@36008.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@36008.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@36008.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@36008.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@36008.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@36017.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@36017.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@36017.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@36017.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@36017.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@36026.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@36026.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@36026.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@36026.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@36026.4]
  wire  b229; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 62:18:@33238.4]
  wire  b230; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 63:18:@33239.4]
  wire  _T_205; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 67:30:@33241.4]
  wire  _T_206; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 67:37:@33242.4]
  wire  _T_210; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 69:76:@33247.4]
  wire  _T_211; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 69:62:@33248.4]
  wire  _T_213; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 69:101:@33249.4]
  wire [31:0] b227_number; // @[Math.scala 723:22:@33223.4 Math.scala 724:14:@33224.4]
  wire [31:0] _T_242; // @[Math.scala 406:49:@33376.4]
  wire [31:0] _T_244; // @[Math.scala 406:56:@33378.4]
  wire [31:0] _T_245; // @[Math.scala 406:56:@33379.4]
  wire [31:0] x410_number; // @[implicits.scala 133:21:@33380.4]
  wire [31:0] _T_255; // @[Math.scala 406:49:@33389.4]
  wire [31:0] _T_257; // @[Math.scala 406:56:@33391.4]
  wire [31:0] _T_258; // @[Math.scala 406:56:@33392.4]
  wire [31:0] b228_number; // @[Math.scala 723:22:@33235.4 Math.scala 724:14:@33236.4]
  wire  _T_262; // @[FixedPoint.scala 50:25:@33398.4]
  wire [15:0] _T_266; // @[Bitwise.scala 72:12:@33400.4]
  wire [15:0] _T_267; // @[FixedPoint.scala 18:52:@33401.4]
  wire  _T_273; // @[Math.scala 451:55:@33403.4]
  wire [15:0] _T_274; // @[FixedPoint.scala 18:52:@33404.4]
  wire  _T_280; // @[Math.scala 451:110:@33406.4]
  wire  _T_281; // @[Math.scala 451:94:@33407.4]
  wire [31:0] _T_283; // @[Cat.scala 30:58:@33409.4]
  wire [31:0] _T_293; // @[Math.scala 406:49:@33417.4]
  wire [31:0] _T_295; // @[Math.scala 406:56:@33419.4]
  wire [31:0] _T_296; // @[Math.scala 406:56:@33420.4]
  wire [31:0] x414_sum_number; // @[Math.scala 154:22:@33431.4 Math.scala 155:14:@33432.4]
  wire  _T_303; // @[FixedPoint.scala 50:25:@33436.4]
  wire [7:0] _T_307; // @[Bitwise.scala 72:12:@33438.4]
  wire [23:0] _T_308; // @[FixedPoint.scala 18:52:@33439.4]
  wire  _T_314; // @[Math.scala 451:55:@33441.4]
  wire [7:0] _T_315; // @[FixedPoint.scala 18:52:@33442.4]
  wire  _T_321; // @[Math.scala 451:110:@33444.4]
  wire  _T_322; // @[Math.scala 451:94:@33445.4]
  wire [31:0] _T_324; // @[Cat.scala 30:58:@33447.4]
  wire [31:0] _T_334; // @[Math.scala 406:49:@33455.4]
  wire [31:0] _T_336; // @[Math.scala 406:56:@33457.4]
  wire [31:0] _T_337; // @[Math.scala 406:56:@33458.4]
  wire [31:0] x417_sum_number; // @[Math.scala 154:22:@33469.4 Math.scala 155:14:@33470.4]
  wire  _T_344; // @[FixedPoint.scala 50:25:@33474.4]
  wire [3:0] _T_348; // @[Bitwise.scala 72:12:@33476.4]
  wire [27:0] _T_349; // @[FixedPoint.scala 18:52:@33477.4]
  wire  _T_355; // @[Math.scala 451:55:@33479.4]
  wire [3:0] _T_356; // @[FixedPoint.scala 18:52:@33480.4]
  wire  _T_362; // @[Math.scala 451:110:@33482.4]
  wire  _T_363; // @[Math.scala 451:94:@33483.4]
  wire [31:0] _T_365; // @[Cat.scala 30:58:@33485.4]
  wire [31:0] _T_375; // @[Math.scala 406:49:@33493.4]
  wire [31:0] _T_377; // @[Math.scala 406:56:@33495.4]
  wire [31:0] _T_378; // @[Math.scala 406:56:@33496.4]
  wire [31:0] x420_sum_number; // @[Math.scala 154:22:@33507.4 Math.scala 155:14:@33508.4]
  wire  _T_385; // @[FixedPoint.scala 50:25:@33512.4]
  wire [1:0] _T_389; // @[Bitwise.scala 72:12:@33514.4]
  wire [29:0] _T_390; // @[FixedPoint.scala 18:52:@33515.4]
  wire  _T_396; // @[Math.scala 451:55:@33517.4]
  wire [1:0] _T_397; // @[FixedPoint.scala 18:52:@33518.4]
  wire  _T_403; // @[Math.scala 451:110:@33520.4]
  wire  _T_404; // @[Math.scala 451:94:@33521.4]
  wire [31:0] _T_406; // @[Cat.scala 30:58:@33523.4]
  wire [31:0] _T_416; // @[Math.scala 406:49:@33531.4]
  wire [31:0] _T_418; // @[Math.scala 406:56:@33533.4]
  wire [31:0] _T_419; // @[Math.scala 406:56:@33534.4]
  wire [31:0] x423_sum_number; // @[Math.scala 154:22:@33545.4 Math.scala 155:14:@33546.4]
  wire  _T_426; // @[FixedPoint.scala 50:25:@33550.4]
  wire [1:0] _T_430; // @[Bitwise.scala 72:12:@33552.4]
  wire [29:0] _T_431; // @[FixedPoint.scala 18:52:@33553.4]
  wire  _T_437; // @[Math.scala 451:55:@33555.4]
  wire [1:0] _T_438; // @[FixedPoint.scala 18:52:@33556.4]
  wire  _T_444; // @[Math.scala 451:110:@33558.4]
  wire  _T_445; // @[Math.scala 451:94:@33559.4]
  wire [31:0] _T_449; // @[package.scala 96:25:@33567.4 package.scala 96:25:@33568.4]
  wire [31:0] _T_459; // @[Math.scala 406:49:@33576.4]
  wire [31:0] _T_461; // @[Math.scala 406:56:@33578.4]
  wire [31:0] _T_462; // @[Math.scala 406:56:@33579.4]
  wire [31:0] _T_466; // @[package.scala 96:25:@33587.4]
  wire [31:0] x426_sum_number; // @[Math.scala 154:22:@33599.4 Math.scala 155:14:@33600.4]
  wire  _T_473; // @[FixedPoint.scala 50:25:@33604.4]
  wire [1:0] _T_477; // @[Bitwise.scala 72:12:@33606.4]
  wire [29:0] _T_478; // @[FixedPoint.scala 18:52:@33607.4]
  wire  _T_484; // @[Math.scala 451:55:@33609.4]
  wire [1:0] _T_485; // @[FixedPoint.scala 18:52:@33610.4]
  wire  _T_491; // @[Math.scala 451:110:@33612.4]
  wire  _T_492; // @[Math.scala 451:94:@33613.4]
  wire [31:0] _T_494; // @[Cat.scala 30:58:@33615.4]
  wire [31:0] _T_504; // @[Math.scala 406:49:@33623.4]
  wire [31:0] _T_506; // @[Math.scala 406:56:@33625.4]
  wire [31:0] _T_507; // @[Math.scala 406:56:@33626.4]
  wire [31:0] x429_sum_number; // @[Math.scala 154:22:@33637.4 Math.scala 155:14:@33638.4]
  wire [31:0] _T_517; // @[Math.scala 476:37:@33643.4]
  wire  x498_x430_D1; // @[package.scala 96:25:@33681.4 package.scala 96:25:@33682.4]
  wire [31:0] x499_x429_sum_D1_number; // @[package.scala 96:25:@33690.4 package.scala 96:25:@33691.4]
  wire [31:0] x432_sub_number; // @[Math.scala 195:22:@33663.4 Math.scala 196:14:@33664.4]
  wire  _T_548; // @[FixedPoint.scala 50:25:@33698.4]
  wire [1:0] _T_552; // @[Bitwise.scala 72:12:@33700.4]
  wire [29:0] _T_553; // @[FixedPoint.scala 18:52:@33701.4]
  wire  _T_559; // @[Math.scala 451:55:@33703.4]
  wire [1:0] _T_560; // @[FixedPoint.scala 18:52:@33704.4]
  wire  _T_566; // @[Math.scala 451:110:@33706.4]
  wire  _T_567; // @[Math.scala 451:94:@33707.4]
  wire [31:0] _T_569; // @[Cat.scala 30:58:@33709.4]
  wire [31:0] x240_1_number; // @[Math.scala 454:20:@33710.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@33715.4]
  wire [40:0] _T_574; // @[Math.scala 461:32:@33715.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@33720.4]
  wire [38:0] _T_577; // @[Math.scala 461:32:@33720.4]
  wire  _T_610; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:101:@33809.4]
  wire  _T_614; // @[package.scala 96:25:@33817.4 package.scala 96:25:@33818.4]
  wire  _T_616; // @[implicits.scala 55:10:@33819.4]
  wire  _T_617; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:118:@33820.4]
  wire  _T_619; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:207:@33822.4]
  wire  _T_620; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:226:@33823.4]
  wire  x502_b229_D21; // @[package.scala 96:25:@33779.4 package.scala 96:25:@33780.4]
  wire  _T_621; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:252:@33824.4]
  wire  x504_b230_D21; // @[package.scala 96:25:@33797.4 package.scala 96:25:@33798.4]
  wire [31:0] x506_b227_D23_number; // @[package.scala 96:25:@33838.4 package.scala 96:25:@33839.4]
  wire [31:0] _T_633; // @[Math.scala 476:37:@33846.4]
  wire [31:0] x507_b228_D23_number; // @[package.scala 96:25:@33863.4 package.scala 96:25:@33864.4]
  wire [31:0] _T_646; // @[Math.scala 476:37:@33869.4]
  wire  x246; // @[package.scala 96:25:@33854.4 package.scala 96:25:@33855.4]
  wire  x247; // @[package.scala 96:25:@33877.4 package.scala 96:25:@33878.4]
  wire  x248; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 183:24:@33881.4]
  wire  _T_684; // @[package.scala 96:25:@33949.4 package.scala 96:25:@33950.4]
  wire  _T_686; // @[implicits.scala 55:10:@33951.4]
  wire  _T_687; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 202:194:@33952.4]
  wire  x508_x249_D21; // @[package.scala 96:25:@33892.4 package.scala 96:25:@33893.4]
  wire  _T_688; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 202:283:@33953.4]
  wire  x511_b229_D45; // @[package.scala 96:25:@33919.4 package.scala 96:25:@33920.4]
  wire  _T_689; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 202:291:@33954.4]
  wire  x512_b230_D45; // @[package.scala 96:25:@33928.4 package.scala 96:25:@33929.4]
  wire [31:0] x252_rdcol_number; // @[Math.scala 195:22:@33973.4 Math.scala 196:14:@33974.4]
  wire [31:0] _T_704; // @[Math.scala 476:37:@33979.4]
  wire  x514_x246_D1; // @[package.scala 96:25:@33996.4 package.scala 96:25:@33997.4]
  wire  x253; // @[package.scala 96:25:@33987.4 package.scala 96:25:@33988.4]
  wire  x254; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 212:24:@34000.4]
  wire  _T_718; // @[FixedPoint.scala 50:25:@34007.4]
  wire [15:0] _T_722; // @[Bitwise.scala 72:12:@34009.4]
  wire [15:0] _T_723; // @[FixedPoint.scala 18:52:@34010.4]
  wire  _T_729; // @[Math.scala 451:55:@34012.4]
  wire [15:0] _T_730; // @[FixedPoint.scala 18:52:@34013.4]
  wire  _T_736; // @[Math.scala 451:110:@34015.4]
  wire  _T_737; // @[Math.scala 451:94:@34016.4]
  wire [31:0] _T_739; // @[Cat.scala 30:58:@34018.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@34028.4]
  wire [31:0] _T_752; // @[Math.scala 406:56:@34029.4]
  wire [31:0] x439_sum_number; // @[Math.scala 154:22:@34040.4 Math.scala 155:14:@34041.4]
  wire  _T_759; // @[FixedPoint.scala 50:25:@34045.4]
  wire [7:0] _T_763; // @[Bitwise.scala 72:12:@34047.4]
  wire [23:0] _T_764; // @[FixedPoint.scala 18:52:@34048.4]
  wire  _T_770; // @[Math.scala 451:55:@34050.4]
  wire [7:0] _T_771; // @[FixedPoint.scala 18:52:@34051.4]
  wire  _T_777; // @[Math.scala 451:110:@34053.4]
  wire  _T_778; // @[Math.scala 451:94:@34054.4]
  wire [31:0] _T_782; // @[package.scala 96:25:@34062.4 package.scala 96:25:@34063.4]
  wire [31:0] _T_792; // @[Math.scala 406:49:@34071.4]
  wire [31:0] _T_794; // @[Math.scala 406:56:@34073.4]
  wire [31:0] _T_795; // @[Math.scala 406:56:@34074.4]
  wire [31:0] _T_799; // @[package.scala 96:25:@34082.4]
  wire [31:0] x442_sum_number; // @[Math.scala 154:22:@34094.4 Math.scala 155:14:@34095.4]
  wire  _T_806; // @[FixedPoint.scala 50:25:@34099.4]
  wire [3:0] _T_810; // @[Bitwise.scala 72:12:@34101.4]
  wire [27:0] _T_811; // @[FixedPoint.scala 18:52:@34102.4]
  wire  _T_817; // @[Math.scala 451:55:@34104.4]
  wire [3:0] _T_818; // @[FixedPoint.scala 18:52:@34105.4]
  wire  _T_824; // @[Math.scala 451:110:@34107.4]
  wire  _T_825; // @[Math.scala 451:94:@34108.4]
  wire [31:0] _T_827; // @[Cat.scala 30:58:@34110.4]
  wire [31:0] _T_837; // @[Math.scala 406:49:@34118.4]
  wire [31:0] _T_839; // @[Math.scala 406:56:@34120.4]
  wire [31:0] _T_840; // @[Math.scala 406:56:@34121.4]
  wire [31:0] x445_sum_number; // @[Math.scala 154:22:@34132.4 Math.scala 155:14:@34133.4]
  wire  _T_847; // @[FixedPoint.scala 50:25:@34137.4]
  wire [1:0] _T_851; // @[Bitwise.scala 72:12:@34139.4]
  wire [29:0] _T_852; // @[FixedPoint.scala 18:52:@34140.4]
  wire  _T_858; // @[Math.scala 451:55:@34142.4]
  wire [1:0] _T_859; // @[FixedPoint.scala 18:52:@34143.4]
  wire  _T_865; // @[Math.scala 451:110:@34145.4]
  wire  _T_866; // @[Math.scala 451:94:@34146.4]
  wire [31:0] _T_868; // @[Cat.scala 30:58:@34148.4]
  wire [31:0] _T_878; // @[Math.scala 406:49:@34156.4]
  wire [31:0] _T_880; // @[Math.scala 406:56:@34158.4]
  wire [31:0] _T_881; // @[Math.scala 406:56:@34159.4]
  wire [31:0] x448_sum_number; // @[Math.scala 154:22:@34170.4 Math.scala 155:14:@34171.4]
  wire  _T_888; // @[FixedPoint.scala 50:25:@34175.4]
  wire [1:0] _T_892; // @[Bitwise.scala 72:12:@34177.4]
  wire [29:0] _T_893; // @[FixedPoint.scala 18:52:@34178.4]
  wire  _T_899; // @[Math.scala 451:55:@34180.4]
  wire [1:0] _T_900; // @[FixedPoint.scala 18:52:@34181.4]
  wire  _T_906; // @[Math.scala 451:110:@34183.4]
  wire  _T_907; // @[Math.scala 451:94:@34184.4]
  wire [31:0] _T_909; // @[Cat.scala 30:58:@34186.4]
  wire [31:0] _T_919; // @[Math.scala 406:49:@34194.4]
  wire [31:0] _T_921; // @[Math.scala 406:56:@34196.4]
  wire [31:0] _T_922; // @[Math.scala 406:56:@34197.4]
  wire [31:0] x451_sum_number; // @[Math.scala 154:22:@34208.4 Math.scala 155:14:@34209.4]
  wire  _T_929; // @[FixedPoint.scala 50:25:@34213.4]
  wire [1:0] _T_933; // @[Bitwise.scala 72:12:@34215.4]
  wire [29:0] _T_934; // @[FixedPoint.scala 18:52:@34216.4]
  wire  _T_940; // @[Math.scala 451:55:@34218.4]
  wire [1:0] _T_941; // @[FixedPoint.scala 18:52:@34219.4]
  wire  _T_947; // @[Math.scala 451:110:@34221.4]
  wire  _T_948; // @[Math.scala 451:94:@34222.4]
  wire [31:0] _T_950; // @[Cat.scala 30:58:@34224.4]
  wire [31:0] _T_960; // @[Math.scala 406:49:@34232.4]
  wire [31:0] _T_962; // @[Math.scala 406:56:@34234.4]
  wire [31:0] _T_963; // @[Math.scala 406:56:@34235.4]
  wire [31:0] x454_sum_number; // @[Math.scala 154:22:@34246.4 Math.scala 155:14:@34247.4]
  wire [31:0] _T_973; // @[Math.scala 476:37:@34252.4]
  wire  x455; // @[package.scala 96:25:@34260.4 package.scala 96:25:@34261.4]
  wire [31:0] x515_x454_sum_D1_number; // @[package.scala 96:25:@34295.4 package.scala 96:25:@34296.4]
  wire [31:0] x457_sub_number; // @[Math.scala 195:22:@34286.4 Math.scala 196:14:@34287.4]
  wire  _T_1030; // @[package.scala 96:25:@34359.4 package.scala 96:25:@34360.4]
  wire  _T_1032; // @[implicits.scala 55:10:@34361.4]
  wire  _T_1033; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 275:194:@34362.4]
  wire  x517_x255_D20; // @[package.scala 96:25:@34338.4 package.scala 96:25:@34339.4]
  wire  _T_1034; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 275:283:@34363.4]
  wire  _T_1035; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 275:291:@34364.4]
  wire [31:0] x261_rdcol_number; // @[Math.scala 195:22:@34383.4 Math.scala 196:14:@34384.4]
  wire [31:0] _T_1052; // @[Math.scala 476:37:@34391.4]
  wire  x262; // @[package.scala 96:25:@34399.4 package.scala 96:25:@34400.4]
  wire  x263; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 291:59:@34403.4]
  wire  _T_1063; // @[FixedPoint.scala 50:25:@34410.4]
  wire [15:0] _T_1067; // @[Bitwise.scala 72:12:@34412.4]
  wire [15:0] _T_1068; // @[FixedPoint.scala 18:52:@34413.4]
  wire  _T_1074; // @[Math.scala 451:55:@34415.4]
  wire [15:0] _T_1075; // @[FixedPoint.scala 18:52:@34416.4]
  wire  _T_1081; // @[Math.scala 451:110:@34418.4]
  wire  _T_1082; // @[Math.scala 451:94:@34419.4]
  wire [31:0] _T_1084; // @[Cat.scala 30:58:@34421.4]
  wire [31:0] _T_1096; // @[Math.scala 406:56:@34431.4]
  wire [31:0] _T_1097; // @[Math.scala 406:56:@34432.4]
  wire [31:0] x461_sum_number; // @[Math.scala 154:22:@34443.4 Math.scala 155:14:@34444.4]
  wire  _T_1104; // @[FixedPoint.scala 50:25:@34448.4]
  wire [7:0] _T_1108; // @[Bitwise.scala 72:12:@34450.4]
  wire [23:0] _T_1109; // @[FixedPoint.scala 18:52:@34451.4]
  wire  _T_1115; // @[Math.scala 451:55:@34453.4]
  wire [7:0] _T_1116; // @[FixedPoint.scala 18:52:@34454.4]
  wire  _T_1122; // @[Math.scala 451:110:@34456.4]
  wire  _T_1123; // @[Math.scala 451:94:@34457.4]
  wire [31:0] _T_1127; // @[package.scala 96:25:@34465.4 package.scala 96:25:@34466.4]
  wire [31:0] _T_1137; // @[Math.scala 406:49:@34474.4]
  wire [31:0] _T_1139; // @[Math.scala 406:56:@34476.4]
  wire [31:0] _T_1140; // @[Math.scala 406:56:@34477.4]
  wire [31:0] _T_1144; // @[package.scala 96:25:@34485.4]
  wire [31:0] x464_sum_number; // @[Math.scala 154:22:@34497.4 Math.scala 155:14:@34498.4]
  wire  _T_1151; // @[FixedPoint.scala 50:25:@34502.4]
  wire [3:0] _T_1155; // @[Bitwise.scala 72:12:@34504.4]
  wire [27:0] _T_1156; // @[FixedPoint.scala 18:52:@34505.4]
  wire  _T_1162; // @[Math.scala 451:55:@34507.4]
  wire [3:0] _T_1163; // @[FixedPoint.scala 18:52:@34508.4]
  wire  _T_1169; // @[Math.scala 451:110:@34510.4]
  wire  _T_1170; // @[Math.scala 451:94:@34511.4]
  wire [31:0] _T_1172; // @[Cat.scala 30:58:@34513.4]
  wire [31:0] _T_1182; // @[Math.scala 406:49:@34521.4]
  wire [31:0] _T_1184; // @[Math.scala 406:56:@34523.4]
  wire [31:0] _T_1185; // @[Math.scala 406:56:@34524.4]
  wire [31:0] x467_sum_number; // @[Math.scala 154:22:@34535.4 Math.scala 155:14:@34536.4]
  wire  _T_1192; // @[FixedPoint.scala 50:25:@34540.4]
  wire [1:0] _T_1196; // @[Bitwise.scala 72:12:@34542.4]
  wire [29:0] _T_1197; // @[FixedPoint.scala 18:52:@34543.4]
  wire  _T_1203; // @[Math.scala 451:55:@34545.4]
  wire [1:0] _T_1204; // @[FixedPoint.scala 18:52:@34546.4]
  wire  _T_1210; // @[Math.scala 451:110:@34548.4]
  wire  _T_1211; // @[Math.scala 451:94:@34549.4]
  wire [31:0] _T_1213; // @[Cat.scala 30:58:@34551.4]
  wire [31:0] _T_1223; // @[Math.scala 406:49:@34559.4]
  wire [31:0] _T_1225; // @[Math.scala 406:56:@34561.4]
  wire [31:0] _T_1226; // @[Math.scala 406:56:@34562.4]
  wire [31:0] x470_sum_number; // @[Math.scala 154:22:@34573.4 Math.scala 155:14:@34574.4]
  wire  _T_1233; // @[FixedPoint.scala 50:25:@34578.4]
  wire [1:0] _T_1237; // @[Bitwise.scala 72:12:@34580.4]
  wire [29:0] _T_1238; // @[FixedPoint.scala 18:52:@34581.4]
  wire  _T_1244; // @[Math.scala 451:55:@34583.4]
  wire [1:0] _T_1245; // @[FixedPoint.scala 18:52:@34584.4]
  wire  _T_1251; // @[Math.scala 451:110:@34586.4]
  wire  _T_1252; // @[Math.scala 451:94:@34587.4]
  wire [31:0] _T_1254; // @[Cat.scala 30:58:@34589.4]
  wire [31:0] _T_1264; // @[Math.scala 406:49:@34597.4]
  wire [31:0] _T_1266; // @[Math.scala 406:56:@34599.4]
  wire [31:0] _T_1267; // @[Math.scala 406:56:@34600.4]
  wire [31:0] x473_sum_number; // @[Math.scala 154:22:@34611.4 Math.scala 155:14:@34612.4]
  wire  _T_1274; // @[FixedPoint.scala 50:25:@34616.4]
  wire [1:0] _T_1278; // @[Bitwise.scala 72:12:@34618.4]
  wire [29:0] _T_1279; // @[FixedPoint.scala 18:52:@34619.4]
  wire  _T_1285; // @[Math.scala 451:55:@34621.4]
  wire [1:0] _T_1286; // @[FixedPoint.scala 18:52:@34622.4]
  wire  _T_1292; // @[Math.scala 451:110:@34624.4]
  wire  _T_1293; // @[Math.scala 451:94:@34625.4]
  wire [31:0] _T_1295; // @[Cat.scala 30:58:@34627.4]
  wire [31:0] _T_1305; // @[Math.scala 406:49:@34635.4]
  wire [31:0] _T_1307; // @[Math.scala 406:56:@34637.4]
  wire [31:0] _T_1308; // @[Math.scala 406:56:@34638.4]
  wire [31:0] x476_sum_number; // @[Math.scala 154:22:@34649.4 Math.scala 155:14:@34650.4]
  wire [31:0] _T_1318; // @[Math.scala 476:37:@34655.4]
  wire  x477; // @[package.scala 96:25:@34663.4 package.scala 96:25:@34664.4]
  wire [31:0] x519_x476_sum_D1_number; // @[package.scala 96:25:@34698.4 package.scala 96:25:@34699.4]
  wire [31:0] x479_sub_number; // @[Math.scala 195:22:@34689.4 Math.scala 196:14:@34690.4]
  wire  _T_1372; // @[package.scala 96:25:@34753.4 package.scala 96:25:@34754.4]
  wire  _T_1374; // @[implicits.scala 55:10:@34755.4]
  wire  _T_1375; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 352:194:@34756.4]
  wire  x521_x264_D20; // @[package.scala 96:25:@34741.4 package.scala 96:25:@34742.4]
  wire  _T_1376; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 352:283:@34757.4]
  wire  _T_1377; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 352:291:@34758.4]
  wire [31:0] x270_rdrow_number; // @[Math.scala 195:22:@34777.4 Math.scala 196:14:@34778.4]
  wire [31:0] _T_1394; // @[Math.scala 406:49:@34784.4]
  wire [31:0] _T_1396; // @[Math.scala 406:56:@34786.4]
  wire [31:0] _T_1397; // @[Math.scala 406:56:@34787.4]
  wire [31:0] x481_number; // @[implicits.scala 133:21:@34788.4]
  wire  x272; // @[package.scala 96:25:@34802.4 package.scala 96:25:@34803.4]
  wire  x522_x247_D1; // @[package.scala 96:25:@34811.4 package.scala 96:25:@34812.4]
  wire  x273; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 364:24:@34815.4]
  wire [31:0] _T_1423; // @[Math.scala 406:49:@34824.4]
  wire [31:0] _T_1425; // @[Math.scala 406:56:@34826.4]
  wire [31:0] _T_1426; // @[Math.scala 406:56:@34827.4]
  wire [31:0] _T_1430; // @[package.scala 96:25:@34835.4]
  wire  _T_1434; // @[FixedPoint.scala 50:25:@34842.4]
  wire [1:0] _T_1438; // @[Bitwise.scala 72:12:@34844.4]
  wire [29:0] _T_1439; // @[FixedPoint.scala 18:52:@34845.4]
  wire  _T_1445; // @[Math.scala 451:55:@34847.4]
  wire [1:0] _T_1446; // @[FixedPoint.scala 18:52:@34848.4]
  wire  _T_1452; // @[Math.scala 451:110:@34850.4]
  wire  _T_1453; // @[Math.scala 451:94:@34851.4]
  wire [31:0] _T_1457; // @[package.scala 96:25:@34859.4 package.scala 96:25:@34860.4]
  wire [31:0] x276_1_number; // @[Math.scala 454:20:@34861.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@34866.4]
  wire [40:0] _T_1462; // @[Math.scala 461:32:@34866.4]
  wire [38:0] _GEN_3; // @[Math.scala 461:32:@34871.4]
  wire [38:0] _T_1465; // @[Math.scala 461:32:@34871.4]
  wire  _T_1498; // @[package.scala 96:25:@34948.4 package.scala 96:25:@34949.4]
  wire  _T_1500; // @[implicits.scala 55:10:@34950.4]
  wire  _T_1501; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 399:194:@34951.4]
  wire  x525_x274_D20; // @[package.scala 96:25:@34918.4 package.scala 96:25:@34919.4]
  wire  _T_1502; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 399:283:@34952.4]
  wire  _T_1503; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 399:326:@34953.4]
  wire  x281; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 403:59:@34964.4]
  wire  _T_1532; // @[package.scala 96:25:@35008.4 package.scala 96:25:@35009.4]
  wire  _T_1534; // @[implicits.scala 55:10:@35010.4]
  wire  _T_1535; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 418:194:@35011.4]
  wire  x529_x282_D20; // @[package.scala 96:25:@34996.4 package.scala 96:25:@34997.4]
  wire  _T_1536; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 418:283:@35012.4]
  wire  _T_1537; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 418:291:@35013.4]
  wire  x286; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 422:59:@35024.4]
  wire  _T_1561; // @[package.scala 96:25:@35057.4 package.scala 96:25:@35058.4]
  wire  _T_1563; // @[implicits.scala 55:10:@35059.4]
  wire  _T_1564; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 433:194:@35060.4]
  wire  x530_x287_D20; // @[package.scala 96:25:@35045.4 package.scala 96:25:@35046.4]
  wire  _T_1565; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 433:283:@35061.4]
  wire  _T_1566; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 433:291:@35062.4]
  wire [31:0] x291_rdrow_number; // @[Math.scala 195:22:@35081.4 Math.scala 196:14:@35082.4]
  wire [31:0] _T_1583; // @[Math.scala 406:49:@35088.4]
  wire [31:0] _T_1585; // @[Math.scala 406:56:@35090.4]
  wire [31:0] _T_1586; // @[Math.scala 406:56:@35091.4]
  wire [31:0] x486_number; // @[implicits.scala 133:21:@35092.4]
  wire  x293; // @[package.scala 96:25:@35106.4 package.scala 96:25:@35107.4]
  wire  x294; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 443:24:@35110.4]
  wire [31:0] _T_1609; // @[Math.scala 406:49:@35119.4]
  wire [31:0] _T_1611; // @[Math.scala 406:56:@35121.4]
  wire [31:0] _T_1612; // @[Math.scala 406:56:@35122.4]
  wire [31:0] _T_1616; // @[package.scala 96:25:@35130.4]
  wire  _T_1620; // @[FixedPoint.scala 50:25:@35137.4]
  wire [1:0] _T_1624; // @[Bitwise.scala 72:12:@35139.4]
  wire [29:0] _T_1625; // @[FixedPoint.scala 18:52:@35140.4]
  wire  _T_1631; // @[Math.scala 451:55:@35142.4]
  wire [1:0] _T_1632; // @[FixedPoint.scala 18:52:@35143.4]
  wire  _T_1638; // @[Math.scala 451:110:@35145.4]
  wire  _T_1639; // @[Math.scala 451:94:@35146.4]
  wire [31:0] _T_1643; // @[package.scala 96:25:@35154.4 package.scala 96:25:@35155.4]
  wire [31:0] x297_1_number; // @[Math.scala 454:20:@35156.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@35161.4]
  wire [40:0] _T_1648; // @[Math.scala 461:32:@35161.4]
  wire [38:0] _GEN_5; // @[Math.scala 461:32:@35166.4]
  wire [38:0] _T_1651; // @[Math.scala 461:32:@35166.4]
  wire  _T_1681; // @[package.scala 96:25:@35234.4 package.scala 96:25:@35235.4]
  wire  _T_1683; // @[implicits.scala 55:10:@35236.4]
  wire  _T_1684; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 470:194:@35237.4]
  wire  x534_x295_D20; // @[package.scala 96:25:@35222.4 package.scala 96:25:@35223.4]
  wire  _T_1685; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 470:283:@35238.4]
  wire  _T_1686; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 470:291:@35239.4]
  wire  x302; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 474:24:@35250.4]
  wire  _T_1713; // @[package.scala 96:25:@35292.4 package.scala 96:25:@35293.4]
  wire  _T_1715; // @[implicits.scala 55:10:@35294.4]
  wire  _T_1716; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 487:194:@35295.4]
  wire  x536_x303_D20; // @[package.scala 96:25:@35280.4 package.scala 96:25:@35281.4]
  wire  _T_1717; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 487:283:@35296.4]
  wire  _T_1718; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 487:291:@35297.4]
  wire  x307; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 491:24:@35308.4]
  wire  _T_1742; // @[package.scala 96:25:@35341.4 package.scala 96:25:@35342.4]
  wire  _T_1744; // @[implicits.scala 55:10:@35343.4]
  wire  _T_1745; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 502:194:@35344.4]
  wire  x537_x308_D20; // @[package.scala 96:25:@35329.4 package.scala 96:25:@35330.4]
  wire  _T_1746; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 502:283:@35345.4]
  wire  _T_1747; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 502:291:@35346.4]
  wire  _T_1878; // @[package.scala 96:25:@35647.4 package.scala 96:25:@35648.4]
  wire  _T_1880; // @[implicits.scala 55:10:@35649.4]
  wire  _T_1881; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:167:@35650.4]
  wire  _T_1883; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:256:@35652.4]
  wire  _T_1884; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:275:@35653.4]
  wire  x541_b229_D64; // @[package.scala 96:25:@35609.4 package.scala 96:25:@35610.4]
  wire  _T_1885; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:301:@35654.4]
  wire  x542_b230_D64; // @[package.scala 96:25:@35618.4 package.scala 96:25:@35619.4]
  wire  _T_1916; // @[package.scala 96:25:@35725.4 package.scala 96:25:@35726.4]
  wire  _T_1918; // @[implicits.scala 55:10:@35727.4]
  wire  _T_1919; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 590:195:@35728.4]
  wire  x545_x249_D41; // @[package.scala 96:25:@35668.4 package.scala 96:25:@35669.4]
  wire  _T_1920; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 590:284:@35729.4]
  wire  x548_b229_D65; // @[package.scala 96:25:@35695.4 package.scala 96:25:@35696.4]
  wire  _T_1921; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 590:292:@35730.4]
  wire  x549_b230_D65; // @[package.scala 96:25:@35704.4 package.scala 96:25:@35705.4]
  wire  _T_1944; // @[package.scala 96:25:@35776.4 package.scala 96:25:@35777.4]
  wire  _T_1946; // @[implicits.scala 55:10:@35778.4]
  wire  _T_1947; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 603:195:@35779.4]
  wire  x551_x255_D40; // @[package.scala 96:25:@35746.4 package.scala 96:25:@35747.4]
  wire  _T_1948; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 603:284:@35780.4]
  wire  _T_1949; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 603:292:@35781.4]
  wire  _T_1972; // @[package.scala 96:25:@35827.4 package.scala 96:25:@35828.4]
  wire  _T_1974; // @[implicits.scala 55:10:@35829.4]
  wire  _T_1975; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 616:195:@35830.4]
  wire  x554_x274_D40; // @[package.scala 96:25:@35797.4 package.scala 96:25:@35798.4]
  wire  _T_1976; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 616:284:@35831.4]
  wire  _T_1977; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 616:292:@35832.4]
  wire  _T_1997; // @[package.scala 96:25:@35869.4 package.scala 96:25:@35870.4]
  wire  _T_1999; // @[implicits.scala 55:10:@35871.4]
  wire  _T_2000; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 627:195:@35872.4]
  wire  x557_x282_D40; // @[package.scala 96:25:@35848.4 package.scala 96:25:@35849.4]
  wire  _T_2001; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 627:284:@35873.4]
  wire  _T_2002; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 627:292:@35874.4]
  wire  _T_2076; // @[package.scala 96:25:@36031.4 package.scala 96:25:@36032.4]
  wire  _T_2078; // @[implicits.scala 55:10:@36033.4]
  wire  x560_b229_D84; // @[package.scala 96:25:@36022.4 package.scala 96:25:@36023.4]
  wire  _T_2079; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 667:117:@36034.4]
  wire  x559_b230_D84; // @[package.scala 96:25:@36013.4 package.scala 96:25:@36014.4]
  wire  _T_2080; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 667:123:@36035.4]
  wire [31:0] x243_sum_number; // @[Math.scala 154:22:@33761.4 Math.scala 155:14:@33762.4]
  wire [31:0] x501_x411_D21_number; // @[package.scala 96:25:@33770.4 package.scala 96:25:@33771.4]
  wire [31:0] x505_x433_D13_number; // @[package.scala 96:25:@33806.4 package.scala 96:25:@33807.4]
  wire [31:0] x509_x411_D45_number; // @[package.scala 96:25:@33901.4 package.scala 96:25:@33902.4]
  wire [31:0] x510_x243_sum_D24_number; // @[package.scala 96:25:@33910.4 package.scala 96:25:@33911.4]
  wire [31:0] x513_x433_D37_number; // @[package.scala 96:25:@33937.4 package.scala 96:25:@33938.4]
  wire [31:0] x258_sum_number; // @[Math.scala 154:22:@34329.4 Math.scala 155:14:@34330.4]
  wire [31:0] x518_x458_D13_number; // @[package.scala 96:25:@34347.4 package.scala 96:25:@34348.4]
  wire [31:0] x267_sum_number; // @[Math.scala 154:22:@34723.4 Math.scala 155:14:@34724.4]
  wire [31:0] x520_x480_D13_number; // @[package.scala 96:25:@34732.4 package.scala 96:25:@34733.4]
  wire [31:0] x526_x278_sum_D1_number; // @[package.scala 96:25:@34927.4 package.scala 96:25:@34928.4]
  wire [31:0] x527_x482_D20_number; // @[package.scala 96:25:@34936.4 package.scala 96:25:@34937.4]
  wire [31:0] x283_sum_number; // @[Math.scala 154:22:@34987.4 Math.scala 155:14:@34988.4]
  wire [31:0] x288_sum_number; // @[Math.scala 154:22:@35036.4 Math.scala 155:14:@35037.4]
  wire [31:0] x532_x299_sum_D1_number; // @[package.scala 96:25:@35204.4 package.scala 96:25:@35205.4]
  wire [31:0] x533_x487_D20_number; // @[package.scala 96:25:@35213.4 package.scala 96:25:@35214.4]
  wire [31:0] x304_sum_number; // @[Math.scala 154:22:@35271.4 Math.scala 155:14:@35272.4]
  wire [31:0] x309_sum_number; // @[Math.scala 154:22:@35320.4 Math.scala 155:14:@35321.4]
  wire [31:0] x539_x411_D64_number; // @[package.scala 96:25:@35591.4 package.scala 96:25:@35592.4]
  wire [31:0] x540_x243_sum_D43_number; // @[package.scala 96:25:@35600.4 package.scala 96:25:@35601.4]
  wire [31:0] x544_x433_D56_number; // @[package.scala 96:25:@35636.4 package.scala 96:25:@35637.4]
  wire [31:0] x546_x411_D65_number; // @[package.scala 96:25:@35677.4 package.scala 96:25:@35678.4]
  wire [31:0] x547_x243_sum_D44_number; // @[package.scala 96:25:@35686.4 package.scala 96:25:@35687.4]
  wire [31:0] x550_x433_D57_number; // @[package.scala 96:25:@35713.4 package.scala 96:25:@35714.4]
  wire [31:0] x552_x458_D33_number; // @[package.scala 96:25:@35755.4 package.scala 96:25:@35756.4]
  wire [31:0] x553_x258_sum_D20_number; // @[package.scala 96:25:@35764.4 package.scala 96:25:@35765.4]
  wire [31:0] x555_x278_sum_D21_number; // @[package.scala 96:25:@35806.4 package.scala 96:25:@35807.4]
  wire [31:0] x556_x482_D40_number; // @[package.scala 96:25:@35815.4 package.scala 96:25:@35816.4]
  wire [31:0] x558_x283_sum_D20_number; // @[package.scala 96:25:@35857.4 package.scala 96:25:@35858.4]
  _ _ ( // @[Math.scala 720:24:@33218.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@33230.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@33253.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x233_lb_0 x233_lb_0 ( // @[m_x233_lb_0.scala 35:17:@33263.4]
    .clock(x233_lb_0_clock),
    .reset(x233_lb_0_reset),
    .io_rPort_8_banks_1(x233_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x233_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x233_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x233_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x233_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x233_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x233_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x233_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x233_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x233_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x233_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x233_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x233_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x233_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x233_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x233_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x233_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x233_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x233_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x233_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x233_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x233_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x233_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x233_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x233_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x233_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x233_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x233_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x233_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x233_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x233_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x233_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x233_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x233_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x233_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x233_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x233_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x233_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x233_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x233_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x233_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x233_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x233_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x233_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x233_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x233_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x233_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x233_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x233_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x233_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x233_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x233_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x233_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x233_lb_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x233_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x233_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x233_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x233_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x233_lb_0_io_wPort_0_en_0)
  );
  x234_lb2_0 x234_lb2_0 ( // @[m_x234_lb2_0.scala 30:17:@33330.4]
    .clock(x234_lb2_0_clock),
    .reset(x234_lb2_0_reset),
    .io_rPort_3_banks_1(x234_lb2_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x234_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x234_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x234_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x234_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x234_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x234_lb2_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x234_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x234_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x234_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x234_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x234_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x234_lb2_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x234_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x234_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x234_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x234_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x234_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x234_lb2_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x234_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x234_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x234_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x234_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x234_lb2_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x234_lb2_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x234_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x234_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x234_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x234_lb2_0_io_wPort_0_en_0)
  );
  x215_sum x414_sum_1 ( // @[Math.scala 150:24:@33425.4]
    .clock(x414_sum_1_clock),
    .reset(x414_sum_1_reset),
    .io_a(x414_sum_1_io_a),
    .io_b(x414_sum_1_io_b),
    .io_flow(x414_sum_1_io_flow),
    .io_result(x414_sum_1_io_result)
  );
  x215_sum x417_sum_1 ( // @[Math.scala 150:24:@33463.4]
    .clock(x417_sum_1_clock),
    .reset(x417_sum_1_reset),
    .io_a(x417_sum_1_io_a),
    .io_b(x417_sum_1_io_b),
    .io_flow(x417_sum_1_io_flow),
    .io_result(x417_sum_1_io_result)
  );
  x215_sum x420_sum_1 ( // @[Math.scala 150:24:@33501.4]
    .clock(x420_sum_1_clock),
    .reset(x420_sum_1_reset),
    .io_a(x420_sum_1_io_a),
    .io_b(x420_sum_1_io_b),
    .io_flow(x420_sum_1_io_flow),
    .io_result(x420_sum_1_io_result)
  );
  x215_sum x423_sum_1 ( // @[Math.scala 150:24:@33539.4]
    .clock(x423_sum_1_clock),
    .reset(x423_sum_1_reset),
    .io_a(x423_sum_1_io_a),
    .io_b(x423_sum_1_io_b),
    .io_flow(x423_sum_1_io_flow),
    .io_result(x423_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@33562.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_2 ( // @[package.scala 93:22:@33580.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x215_sum x426_sum_1 ( // @[Math.scala 150:24:@33593.4]
    .clock(x426_sum_1_clock),
    .reset(x426_sum_1_reset),
    .io_a(x426_sum_1_io_a),
    .io_b(x426_sum_1_io_b),
    .io_flow(x426_sum_1_io_flow),
    .io_result(x426_sum_1_io_result)
  );
  x215_sum x429_sum_1 ( // @[Math.scala 150:24:@33631.4]
    .clock(x429_sum_1_clock),
    .reset(x429_sum_1_reset),
    .io_a(x429_sum_1_io_a),
    .io_b(x429_sum_1_io_b),
    .io_flow(x429_sum_1_io_flow),
    .io_result(x429_sum_1_io_result)
  );
  x408_sub x432_sub_1 ( // @[Math.scala 191:24:@33657.4]
    .clock(x432_sub_1_clock),
    .reset(x432_sub_1_reset),
    .io_a(x432_sub_1_io_a),
    .io_b(x432_sub_1_io_b),
    .io_flow(x432_sub_1_io_flow),
    .io_result(x432_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@33667.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@33676.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_5 ( // @[package.scala 93:22:@33685.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x215_sum x436_sum_1 ( // @[Math.scala 150:24:@33724.4]
    .clock(x436_sum_1_clock),
    .reset(x436_sum_1_reset),
    .io_a(x436_sum_1_io_a),
    .io_b(x436_sum_1_io_b),
    .io_flow(x436_sum_1_io_flow),
    .io_result(x436_sum_1_io_result)
  );
  x242_div x242_div_1 ( // @[Math.scala 327:24:@33736.4]
    .clock(x242_div_1_clock),
    .io_a(x242_div_1_io_a),
    .io_flow(x242_div_1_io_flow),
    .io_result(x242_div_1_io_result)
  );
  RetimeWrapper_243 RetimeWrapper_6 ( // @[package.scala 93:22:@33746.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x215_sum x243_sum_1 ( // @[Math.scala 150:24:@33755.4]
    .clock(x243_sum_1_clock),
    .reset(x243_sum_1_reset),
    .io_a(x243_sum_1_io_a),
    .io_b(x243_sum_1_io_b),
    .io_flow(x243_sum_1_io_flow),
    .io_result(x243_sum_1_io_result)
  );
  RetimeWrapper_245 RetimeWrapper_7 ( // @[package.scala 93:22:@33765.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_8 ( // @[package.scala 93:22:@33774.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_9 ( // @[package.scala 93:22:@33783.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_10 ( // @[package.scala 93:22:@33792.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_11 ( // @[package.scala 93:22:@33801.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_12 ( // @[package.scala 93:22:@33812.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_251 RetimeWrapper_13 ( // @[package.scala 93:22:@33833.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@33849.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_251 RetimeWrapper_15 ( // @[package.scala 93:22:@33858.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@33872.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_17 ( // @[package.scala 93:22:@33887.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_256 RetimeWrapper_18 ( // @[package.scala 93:22:@33896.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_257 RetimeWrapper_19 ( // @[package.scala 93:22:@33905.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_20 ( // @[package.scala 93:22:@33914.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_21 ( // @[package.scala 93:22:@33923.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_260 RetimeWrapper_22 ( // @[package.scala 93:22:@33932.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_23 ( // @[package.scala 93:22:@33944.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  x408_sub x252_rdcol_1 ( // @[Math.scala 191:24:@33967.4]
    .clock(x252_rdcol_1_clock),
    .reset(x252_rdcol_1_reset),
    .io_a(x252_rdcol_1_io_a),
    .io_b(x252_rdcol_1_io_b),
    .io_flow(x252_rdcol_1_io_flow),
    .io_result(x252_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@33982.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@33991.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  x215_sum x439_sum_1 ( // @[Math.scala 150:24:@34034.4]
    .clock(x439_sum_1_clock),
    .reset(x439_sum_1_reset),
    .io_a(x439_sum_1_io_a),
    .io_b(x439_sum_1_io_b),
    .io_flow(x439_sum_1_io_flow),
    .io_result(x439_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_26 ( // @[package.scala 93:22:@34057.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_27 ( // @[package.scala 93:22:@34075.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x215_sum x442_sum_1 ( // @[Math.scala 150:24:@34088.4]
    .clock(x442_sum_1_clock),
    .reset(x442_sum_1_reset),
    .io_a(x442_sum_1_io_a),
    .io_b(x442_sum_1_io_b),
    .io_flow(x442_sum_1_io_flow),
    .io_result(x442_sum_1_io_result)
  );
  x215_sum x445_sum_1 ( // @[Math.scala 150:24:@34126.4]
    .clock(x445_sum_1_clock),
    .reset(x445_sum_1_reset),
    .io_a(x445_sum_1_io_a),
    .io_b(x445_sum_1_io_b),
    .io_flow(x445_sum_1_io_flow),
    .io_result(x445_sum_1_io_result)
  );
  x215_sum x448_sum_1 ( // @[Math.scala 150:24:@34164.4]
    .clock(x448_sum_1_clock),
    .reset(x448_sum_1_reset),
    .io_a(x448_sum_1_io_a),
    .io_b(x448_sum_1_io_b),
    .io_flow(x448_sum_1_io_flow),
    .io_result(x448_sum_1_io_result)
  );
  x215_sum x451_sum_1 ( // @[Math.scala 150:24:@34202.4]
    .clock(x451_sum_1_clock),
    .reset(x451_sum_1_reset),
    .io_a(x451_sum_1_io_a),
    .io_b(x451_sum_1_io_b),
    .io_flow(x451_sum_1_io_flow),
    .io_result(x451_sum_1_io_result)
  );
  x215_sum x454_sum_1 ( // @[Math.scala 150:24:@34240.4]
    .clock(x454_sum_1_clock),
    .reset(x454_sum_1_reset),
    .io_a(x454_sum_1_io_a),
    .io_b(x454_sum_1_io_b),
    .io_flow(x454_sum_1_io_flow),
    .io_result(x454_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@34255.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@34269.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  x408_sub x457_sub_1 ( // @[Math.scala 191:24:@34280.4]
    .clock(x457_sub_1_clock),
    .reset(x457_sub_1_reset),
    .io_a(x457_sub_1_io_a),
    .io_b(x457_sub_1_io_b),
    .io_flow(x457_sub_1_io_flow),
    .io_result(x457_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_30 ( // @[package.scala 93:22:@34290.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x242_div x257_div_1 ( // @[Math.scala 327:24:@34304.4]
    .clock(x257_div_1_clock),
    .io_a(x257_div_1_io_a),
    .io_flow(x257_div_1_io_flow),
    .io_result(x257_div_1_io_result)
  );
  RetimeWrapper_277 RetimeWrapper_31 ( // @[package.scala 93:22:@34314.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x215_sum x258_sum_1 ( // @[Math.scala 150:24:@34323.4]
    .clock(x258_sum_1_clock),
    .reset(x258_sum_1_reset),
    .io_a(x258_sum_1_io_a),
    .io_b(x258_sum_1_io_b),
    .io_flow(x258_sum_1_io_flow),
    .io_result(x258_sum_1_io_result)
  );
  RetimeWrapper_279 RetimeWrapper_32 ( // @[package.scala 93:22:@34333.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_33 ( // @[package.scala 93:22:@34342.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_34 ( // @[package.scala 93:22:@34354.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x408_sub x261_rdcol_1 ( // @[Math.scala 191:24:@34377.4]
    .clock(x261_rdcol_1_clock),
    .reset(x261_rdcol_1_reset),
    .io_a(x261_rdcol_1_io_a),
    .io_b(x261_rdcol_1_io_b),
    .io_flow(x261_rdcol_1_io_flow),
    .io_result(x261_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@34394.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  x215_sum x461_sum_1 ( // @[Math.scala 150:24:@34437.4]
    .clock(x461_sum_1_clock),
    .reset(x461_sum_1_reset),
    .io_a(x461_sum_1_io_a),
    .io_b(x461_sum_1_io_b),
    .io_flow(x461_sum_1_io_flow),
    .io_result(x461_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_36 ( // @[package.scala 93:22:@34460.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_37 ( // @[package.scala 93:22:@34478.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x215_sum x464_sum_1 ( // @[Math.scala 150:24:@34491.4]
    .clock(x464_sum_1_clock),
    .reset(x464_sum_1_reset),
    .io_a(x464_sum_1_io_a),
    .io_b(x464_sum_1_io_b),
    .io_flow(x464_sum_1_io_flow),
    .io_result(x464_sum_1_io_result)
  );
  x215_sum x467_sum_1 ( // @[Math.scala 150:24:@34529.4]
    .clock(x467_sum_1_clock),
    .reset(x467_sum_1_reset),
    .io_a(x467_sum_1_io_a),
    .io_b(x467_sum_1_io_b),
    .io_flow(x467_sum_1_io_flow),
    .io_result(x467_sum_1_io_result)
  );
  x215_sum x470_sum_1 ( // @[Math.scala 150:24:@34567.4]
    .clock(x470_sum_1_clock),
    .reset(x470_sum_1_reset),
    .io_a(x470_sum_1_io_a),
    .io_b(x470_sum_1_io_b),
    .io_flow(x470_sum_1_io_flow),
    .io_result(x470_sum_1_io_result)
  );
  x215_sum x473_sum_1 ( // @[Math.scala 150:24:@34605.4]
    .clock(x473_sum_1_clock),
    .reset(x473_sum_1_reset),
    .io_a(x473_sum_1_io_a),
    .io_b(x473_sum_1_io_b),
    .io_flow(x473_sum_1_io_flow),
    .io_result(x473_sum_1_io_result)
  );
  x215_sum x476_sum_1 ( // @[Math.scala 150:24:@34643.4]
    .clock(x476_sum_1_clock),
    .reset(x476_sum_1_reset),
    .io_a(x476_sum_1_io_a),
    .io_b(x476_sum_1_io_b),
    .io_flow(x476_sum_1_io_flow),
    .io_result(x476_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@34658.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper RetimeWrapper_39 ( // @[package.scala 93:22:@34672.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x408_sub x479_sub_1 ( // @[Math.scala 191:24:@34683.4]
    .clock(x479_sub_1_clock),
    .reset(x479_sub_1_reset),
    .io_a(x479_sub_1_io_a),
    .io_b(x479_sub_1_io_b),
    .io_flow(x479_sub_1_io_flow),
    .io_result(x479_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_40 ( // @[package.scala 93:22:@34693.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x242_div x266_div_1 ( // @[Math.scala 327:24:@34707.4]
    .clock(x266_div_1_clock),
    .io_a(x266_div_1_io_a),
    .io_flow(x266_div_1_io_flow),
    .io_result(x266_div_1_io_result)
  );
  x215_sum x267_sum_1 ( // @[Math.scala 150:24:@34717.4]
    .clock(x267_sum_1_clock),
    .reset(x267_sum_1_reset),
    .io_a(x267_sum_1_io_a),
    .io_b(x267_sum_1_io_b),
    .io_flow(x267_sum_1_io_flow),
    .io_result(x267_sum_1_io_result)
  );
  RetimeWrapper_249 RetimeWrapper_41 ( // @[package.scala 93:22:@34727.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_279 RetimeWrapper_42 ( // @[package.scala 93:22:@34736.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_43 ( // @[package.scala 93:22:@34748.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x408_sub x270_rdrow_1 ( // @[Math.scala 191:24:@34771.4]
    .clock(x270_rdrow_1_clock),
    .reset(x270_rdrow_1_reset),
    .io_a(x270_rdrow_1_io_a),
    .io_b(x270_rdrow_1_io_b),
    .io_flow(x270_rdrow_1_io_flow),
    .io_result(x270_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@34797.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@34806.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_46 ( // @[package.scala 93:22:@34828.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_47 ( // @[package.scala 93:22:@34854.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  x215_sum x485_sum_1 ( // @[Math.scala 150:24:@34875.4]
    .clock(x485_sum_1_clock),
    .reset(x485_sum_1_reset),
    .io_a(x485_sum_1_io_a),
    .io_b(x485_sum_1_io_b),
    .io_flow(x485_sum_1_io_flow),
    .io_result(x485_sum_1_io_result)
  );
  RetimeWrapper_251 RetimeWrapper_48 ( // @[package.scala 93:22:@34885.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_307 RetimeWrapper_49 ( // @[package.scala 93:22:@34894.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  x215_sum x278_sum_1 ( // @[Math.scala 150:24:@34903.4]
    .clock(x278_sum_1_clock),
    .reset(x278_sum_1_reset),
    .io_a(x278_sum_1_io_a),
    .io_b(x278_sum_1_io_b),
    .io_flow(x278_sum_1_io_flow),
    .io_result(x278_sum_1_io_result)
  );
  RetimeWrapper_279 RetimeWrapper_50 ( // @[package.scala 93:22:@34913.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_51 ( // @[package.scala 93:22:@34922.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_52 ( // @[package.scala 93:22:@34931.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_53 ( // @[package.scala 93:22:@34943.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_313 RetimeWrapper_54 ( // @[package.scala 93:22:@34970.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x215_sum x283_sum_1 ( // @[Math.scala 150:24:@34981.4]
    .clock(x283_sum_1_clock),
    .reset(x283_sum_1_reset),
    .io_a(x283_sum_1_io_a),
    .io_b(x283_sum_1_io_b),
    .io_flow(x283_sum_1_io_flow),
    .io_result(x283_sum_1_io_result)
  );
  RetimeWrapper_279 RetimeWrapper_55 ( // @[package.scala 93:22:@34991.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_56 ( // @[package.scala 93:22:@35003.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x215_sum x288_sum_1 ( // @[Math.scala 150:24:@35030.4]
    .clock(x288_sum_1_clock),
    .reset(x288_sum_1_reset),
    .io_a(x288_sum_1_io_a),
    .io_b(x288_sum_1_io_b),
    .io_flow(x288_sum_1_io_flow),
    .io_result(x288_sum_1_io_result)
  );
  RetimeWrapper_279 RetimeWrapper_57 ( // @[package.scala 93:22:@35040.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_58 ( // @[package.scala 93:22:@35052.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x408_sub x291_rdrow_1 ( // @[Math.scala 191:24:@35075.4]
    .clock(x291_rdrow_1_clock),
    .reset(x291_rdrow_1_reset),
    .io_a(x291_rdrow_1_io_a),
    .io_b(x291_rdrow_1_io_b),
    .io_flow(x291_rdrow_1_io_flow),
    .io_result(x291_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_59 ( // @[package.scala 93:22:@35101.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_60 ( // @[package.scala 93:22:@35123.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_61 ( // @[package.scala 93:22:@35149.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x215_sum x490_sum_1 ( // @[Math.scala 150:24:@35170.4]
    .clock(x490_sum_1_clock),
    .reset(x490_sum_1_reset),
    .io_a(x490_sum_1_io_a),
    .io_b(x490_sum_1_io_b),
    .io_flow(x490_sum_1_io_flow),
    .io_result(x490_sum_1_io_result)
  );
  RetimeWrapper_307 RetimeWrapper_62 ( // @[package.scala 93:22:@35180.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x215_sum x299_sum_1 ( // @[Math.scala 150:24:@35189.4]
    .clock(x299_sum_1_clock),
    .reset(x299_sum_1_reset),
    .io_a(x299_sum_1_io_a),
    .io_b(x299_sum_1_io_b),
    .io_flow(x299_sum_1_io_flow),
    .io_result(x299_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_63 ( // @[package.scala 93:22:@35199.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_64 ( // @[package.scala 93:22:@35208.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_279 RetimeWrapper_65 ( // @[package.scala 93:22:@35217.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_66 ( // @[package.scala 93:22:@35229.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_313 RetimeWrapper_67 ( // @[package.scala 93:22:@35256.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x215_sum x304_sum_1 ( // @[Math.scala 150:24:@35265.4]
    .clock(x304_sum_1_clock),
    .reset(x304_sum_1_reset),
    .io_a(x304_sum_1_io_a),
    .io_b(x304_sum_1_io_b),
    .io_flow(x304_sum_1_io_flow),
    .io_result(x304_sum_1_io_result)
  );
  RetimeWrapper_279 RetimeWrapper_68 ( // @[package.scala 93:22:@35275.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_69 ( // @[package.scala 93:22:@35287.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x215_sum x309_sum_1 ( // @[Math.scala 150:24:@35314.4]
    .clock(x309_sum_1_clock),
    .reset(x309_sum_1_reset),
    .io_a(x309_sum_1_io_a),
    .io_b(x309_sum_1_io_b),
    .io_flow(x309_sum_1_io_flow),
    .io_result(x309_sum_1_io_result)
  );
  RetimeWrapper_279 RetimeWrapper_70 ( // @[package.scala 93:22:@35324.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_258 RetimeWrapper_71 ( // @[package.scala 93:22:@35336.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x312 x312_1 ( // @[Math.scala 262:24:@35359.4]
    .clock(x312_1_clock),
    .io_a(x312_1_io_a),
    .io_b(x312_1_io_b),
    .io_flow(x312_1_io_flow),
    .io_result(x312_1_io_result)
  );
  x312 x313_1 ( // @[Math.scala 262:24:@35371.4]
    .clock(x313_1_clock),
    .io_a(x313_1_io_a),
    .io_b(x313_1_io_b),
    .io_flow(x313_1_io_flow),
    .io_result(x313_1_io_result)
  );
  x312 x314_1 ( // @[Math.scala 262:24:@35383.4]
    .clock(x314_1_clock),
    .io_a(x314_1_io_a),
    .io_b(x314_1_io_b),
    .io_flow(x314_1_io_flow),
    .io_result(x314_1_io_result)
  );
  x312 x315_1 ( // @[Math.scala 262:24:@35395.4]
    .clock(x315_1_clock),
    .io_a(x315_1_io_a),
    .io_b(x315_1_io_b),
    .io_flow(x315_1_io_flow),
    .io_result(x315_1_io_result)
  );
  x312 x316_1 ( // @[Math.scala 262:24:@35409.4]
    .clock(x316_1_clock),
    .io_a(x316_1_io_a),
    .io_b(x316_1_io_b),
    .io_flow(x316_1_io_flow),
    .io_result(x316_1_io_result)
  );
  x312 x317_1 ( // @[Math.scala 262:24:@35421.4]
    .clock(x317_1_clock),
    .io_a(x317_1_io_a),
    .io_b(x317_1_io_b),
    .io_flow(x317_1_io_flow),
    .io_result(x317_1_io_result)
  );
  x312 x318_1 ( // @[Math.scala 262:24:@35433.4]
    .clock(x318_1_clock),
    .io_a(x318_1_io_a),
    .io_b(x318_1_io_b),
    .io_flow(x318_1_io_flow),
    .io_result(x318_1_io_result)
  );
  x312 x319_1 ( // @[Math.scala 262:24:@35445.4]
    .clock(x319_1_clock),
    .io_a(x319_1_io_a),
    .io_b(x319_1_io_b),
    .io_flow(x319_1_io_flow),
    .io_result(x319_1_io_result)
  );
  x312 x320_1 ( // @[Math.scala 262:24:@35457.4]
    .clock(x320_1_clock),
    .io_a(x320_1_io_a),
    .io_b(x320_1_io_b),
    .io_flow(x320_1_io_flow),
    .io_result(x320_1_io_result)
  );
  x321_x7 x321_x7_1 ( // @[Math.scala 150:24:@35467.4]
    .clock(x321_x7_1_clock),
    .reset(x321_x7_1_reset),
    .io_a(x321_x7_1_io_a),
    .io_b(x321_x7_1_io_b),
    .io_flow(x321_x7_1_io_flow),
    .io_result(x321_x7_1_io_result)
  );
  x321_x7 x322_x8_1 ( // @[Math.scala 150:24:@35477.4]
    .clock(x322_x8_1_clock),
    .reset(x322_x8_1_reset),
    .io_a(x322_x8_1_io_a),
    .io_b(x322_x8_1_io_b),
    .io_flow(x322_x8_1_io_flow),
    .io_result(x322_x8_1_io_result)
  );
  x321_x7 x323_x7_1 ( // @[Math.scala 150:24:@35487.4]
    .clock(x323_x7_1_clock),
    .reset(x323_x7_1_reset),
    .io_a(x323_x7_1_io_a),
    .io_b(x323_x7_1_io_b),
    .io_flow(x323_x7_1_io_flow),
    .io_result(x323_x7_1_io_result)
  );
  x321_x7 x324_x8_1 ( // @[Math.scala 150:24:@35497.4]
    .clock(x324_x8_1_clock),
    .reset(x324_x8_1_reset),
    .io_a(x324_x8_1_io_a),
    .io_b(x324_x8_1_io_b),
    .io_flow(x324_x8_1_io_flow),
    .io_result(x324_x8_1_io_result)
  );
  x321_x7 x325_x7_1 ( // @[Math.scala 150:24:@35507.4]
    .clock(x325_x7_1_clock),
    .reset(x325_x7_1_reset),
    .io_a(x325_x7_1_io_a),
    .io_b(x325_x7_1_io_b),
    .io_flow(x325_x7_1_io_flow),
    .io_result(x325_x7_1_io_result)
  );
  x321_x7 x326_x8_1 ( // @[Math.scala 150:24:@35517.4]
    .clock(x326_x8_1_clock),
    .reset(x326_x8_1_reset),
    .io_a(x326_x8_1_io_a),
    .io_b(x326_x8_1_io_b),
    .io_flow(x326_x8_1_io_flow),
    .io_result(x326_x8_1_io_result)
  );
  x321_x7 x327_x7_1 ( // @[Math.scala 150:24:@35527.4]
    .clock(x327_x7_1_clock),
    .reset(x327_x7_1_reset),
    .io_a(x327_x7_1_io_a),
    .io_b(x327_x7_1_io_b),
    .io_flow(x327_x7_1_io_flow),
    .io_result(x327_x7_1_io_result)
  );
  RetimeWrapper_345 RetimeWrapper_72 ( // @[package.scala 93:22:@35537.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x321_x7 x328_sum_1 ( // @[Math.scala 150:24:@35546.4]
    .clock(x328_sum_1_clock),
    .reset(x328_sum_1_reset),
    .io_a(x328_sum_1_io_a),
    .io_b(x328_sum_1_io_b),
    .io_flow(x328_sum_1_io_flow),
    .io_result(x328_sum_1_io_result)
  );
  x329 x329_1 ( // @[Math.scala 720:24:@35556.4]
    .io_b(x329_1_io_b),
    .io_result(x329_1_io_result)
  );
  x330_mul x330_mul_1 ( // @[Math.scala 262:24:@35567.4]
    .clock(x330_mul_1_clock),
    .io_a(x330_mul_1_io_a),
    .io_b(x330_mul_1_io_b),
    .io_flow(x330_mul_1_io_flow),
    .io_result(x330_mul_1_io_result)
  );
  x331 x331_1 ( // @[Math.scala 720:24:@35577.4]
    .io_b(x331_1_io_b),
    .io_result(x331_1_io_result)
  );
  RetimeWrapper_347 RetimeWrapper_73 ( // @[package.scala 93:22:@35586.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_277 RetimeWrapper_74 ( // @[package.scala 93:22:@35595.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_75 ( // @[package.scala 93:22:@35604.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_76 ( // @[package.scala 93:22:@35613.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_77 ( // @[package.scala 93:22:@35622.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_78 ( // @[package.scala 93:22:@35631.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_349 RetimeWrapper_79 ( // @[package.scala 93:22:@35642.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_354 RetimeWrapper_80 ( // @[package.scala 93:22:@35663.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_81 ( // @[package.scala 93:22:@35672.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_356 RetimeWrapper_82 ( // @[package.scala 93:22:@35681.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_357 RetimeWrapper_83 ( // @[package.scala 93:22:@35690.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_357 RetimeWrapper_84 ( // @[package.scala 93:22:@35699.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_359 RetimeWrapper_85 ( // @[package.scala 93:22:@35708.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_357 RetimeWrapper_86 ( // @[package.scala 93:22:@35720.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_361 RetimeWrapper_87 ( // @[package.scala 93:22:@35741.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_362 RetimeWrapper_88 ( // @[package.scala 93:22:@35750.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_89 ( // @[package.scala 93:22:@35759.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_357 RetimeWrapper_90 ( // @[package.scala 93:22:@35771.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_361 RetimeWrapper_91 ( // @[package.scala 93:22:@35792.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_245 RetimeWrapper_92 ( // @[package.scala 93:22:@35801.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_367 RetimeWrapper_93 ( // @[package.scala 93:22:@35810.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_357 RetimeWrapper_94 ( // @[package.scala 93:22:@35822.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_361 RetimeWrapper_95 ( // @[package.scala 93:22:@35843.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_96 ( // @[package.scala 93:22:@35852.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_357 RetimeWrapper_97 ( // @[package.scala 93:22:@35864.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  x312 x343_1 ( // @[Math.scala 262:24:@35887.4]
    .clock(x343_1_clock),
    .io_a(x343_1_io_a),
    .io_b(x343_1_io_b),
    .io_flow(x343_1_io_flow),
    .io_result(x343_1_io_result)
  );
  x312 x344_1 ( // @[Math.scala 262:24:@35901.4]
    .clock(x344_1_clock),
    .io_a(x344_1_io_a),
    .io_b(x344_1_io_b),
    .io_flow(x344_1_io_flow),
    .io_result(x344_1_io_result)
  );
  x312 x345_1 ( // @[Math.scala 262:24:@35913.4]
    .clock(x345_1_clock),
    .io_a(x345_1_io_a),
    .io_b(x345_1_io_b),
    .io_flow(x345_1_io_flow),
    .io_result(x345_1_io_result)
  );
  x312 x346_1 ( // @[Math.scala 262:24:@35925.4]
    .clock(x346_1_clock),
    .io_a(x346_1_io_a),
    .io_b(x346_1_io_b),
    .io_flow(x346_1_io_flow),
    .io_result(x346_1_io_result)
  );
  x321_x7 x347_x9_1 ( // @[Math.scala 150:24:@35935.4]
    .clock(x347_x9_1_clock),
    .reset(x347_x9_1_reset),
    .io_a(x347_x9_1_io_a),
    .io_b(x347_x9_1_io_b),
    .io_flow(x347_x9_1_io_flow),
    .io_result(x347_x9_1_io_result)
  );
  x321_x7 x348_x10_1 ( // @[Math.scala 150:24:@35945.4]
    .clock(x348_x10_1_clock),
    .reset(x348_x10_1_reset),
    .io_a(x348_x10_1_io_a),
    .io_b(x348_x10_1_io_b),
    .io_flow(x348_x10_1_io_flow),
    .io_result(x348_x10_1_io_result)
  );
  x321_x7 x349_sum_1 ( // @[Math.scala 150:24:@35955.4]
    .clock(x349_sum_1_clock),
    .reset(x349_sum_1_reset),
    .io_a(x349_sum_1_io_a),
    .io_b(x349_sum_1_io_b),
    .io_flow(x349_sum_1_io_flow),
    .io_result(x349_sum_1_io_result)
  );
  x329 x350_1 ( // @[Math.scala 720:24:@35965.4]
    .io_b(x350_1_io_b),
    .io_result(x350_1_io_result)
  );
  x330_mul x351_mul_1 ( // @[Math.scala 262:24:@35976.4]
    .clock(x351_mul_1_clock),
    .io_a(x351_mul_1_io_a),
    .io_b(x351_mul_1_io_b),
    .io_flow(x351_mul_1_io_flow),
    .io_result(x351_mul_1_io_result)
  );
  x331 x352_1 ( // @[Math.scala 720:24:@35986.4]
    .io_b(x352_1_io_b),
    .io_result(x352_1_io_result)
  );
  RetimeWrapper_345 RetimeWrapper_98 ( // @[package.scala 93:22:@35999.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_376 RetimeWrapper_99 ( // @[package.scala 93:22:@36008.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_376 RetimeWrapper_100 ( // @[package.scala 93:22:@36017.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_376 RetimeWrapper_101 ( // @[package.scala 93:22:@36026.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  assign b229 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 62:18:@33238.4]
  assign b230 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 63:18:@33239.4]
  assign _T_205 = b229 & b230; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 67:30:@33241.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 67:37:@33242.4]
  assign _T_210 = io_in_x201_TID == 8'h0; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 69:76:@33247.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 69:62:@33248.4]
  assign _T_213 = io_in_x201_TDEST == 8'h0; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 69:101:@33249.4]
  assign b227_number = __io_result; // @[Math.scala 723:22:@33223.4 Math.scala 724:14:@33224.4]
  assign _T_242 = $signed(b227_number); // @[Math.scala 406:49:@33376.4]
  assign _T_244 = $signed(_T_242) & $signed(32'sh3); // @[Math.scala 406:56:@33378.4]
  assign _T_245 = $signed(_T_244); // @[Math.scala 406:56:@33379.4]
  assign x410_number = $unsigned(_T_245); // @[implicits.scala 133:21:@33380.4]
  assign _T_255 = $signed(x410_number); // @[Math.scala 406:49:@33389.4]
  assign _T_257 = $signed(_T_255) & $signed(32'sh3); // @[Math.scala 406:56:@33391.4]
  assign _T_258 = $signed(_T_257); // @[Math.scala 406:56:@33392.4]
  assign b228_number = __1_io_result; // @[Math.scala 723:22:@33235.4 Math.scala 724:14:@33236.4]
  assign _T_262 = b228_number[31]; // @[FixedPoint.scala 50:25:@33398.4]
  assign _T_266 = _T_262 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@33400.4]
  assign _T_267 = b228_number[31:16]; // @[FixedPoint.scala 18:52:@33401.4]
  assign _T_273 = _T_267 == 16'hffff; // @[Math.scala 451:55:@33403.4]
  assign _T_274 = b228_number[15:0]; // @[FixedPoint.scala 18:52:@33404.4]
  assign _T_280 = _T_274 != 16'h0; // @[Math.scala 451:110:@33406.4]
  assign _T_281 = _T_273 & _T_280; // @[Math.scala 451:94:@33407.4]
  assign _T_283 = {_T_266,_T_267}; // @[Cat.scala 30:58:@33409.4]
  assign _T_293 = $signed(b228_number); // @[Math.scala 406:49:@33417.4]
  assign _T_295 = $signed(_T_293) & $signed(32'shffff); // @[Math.scala 406:56:@33419.4]
  assign _T_296 = $signed(_T_295); // @[Math.scala 406:56:@33420.4]
  assign x414_sum_number = x414_sum_1_io_result; // @[Math.scala 154:22:@33431.4 Math.scala 155:14:@33432.4]
  assign _T_303 = x414_sum_number[31]; // @[FixedPoint.scala 50:25:@33436.4]
  assign _T_307 = _T_303 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@33438.4]
  assign _T_308 = x414_sum_number[31:8]; // @[FixedPoint.scala 18:52:@33439.4]
  assign _T_314 = _T_308 == 24'hffffff; // @[Math.scala 451:55:@33441.4]
  assign _T_315 = x414_sum_number[7:0]; // @[FixedPoint.scala 18:52:@33442.4]
  assign _T_321 = _T_315 != 8'h0; // @[Math.scala 451:110:@33444.4]
  assign _T_322 = _T_314 & _T_321; // @[Math.scala 451:94:@33445.4]
  assign _T_324 = {_T_307,_T_308}; // @[Cat.scala 30:58:@33447.4]
  assign _T_334 = $signed(x414_sum_number); // @[Math.scala 406:49:@33455.4]
  assign _T_336 = $signed(_T_334) & $signed(32'shff); // @[Math.scala 406:56:@33457.4]
  assign _T_337 = $signed(_T_336); // @[Math.scala 406:56:@33458.4]
  assign x417_sum_number = x417_sum_1_io_result; // @[Math.scala 154:22:@33469.4 Math.scala 155:14:@33470.4]
  assign _T_344 = x417_sum_number[31]; // @[FixedPoint.scala 50:25:@33474.4]
  assign _T_348 = _T_344 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@33476.4]
  assign _T_349 = x417_sum_number[31:4]; // @[FixedPoint.scala 18:52:@33477.4]
  assign _T_355 = _T_349 == 28'hfffffff; // @[Math.scala 451:55:@33479.4]
  assign _T_356 = x417_sum_number[3:0]; // @[FixedPoint.scala 18:52:@33480.4]
  assign _T_362 = _T_356 != 4'h0; // @[Math.scala 451:110:@33482.4]
  assign _T_363 = _T_355 & _T_362; // @[Math.scala 451:94:@33483.4]
  assign _T_365 = {_T_348,_T_349}; // @[Cat.scala 30:58:@33485.4]
  assign _T_375 = $signed(x417_sum_number); // @[Math.scala 406:49:@33493.4]
  assign _T_377 = $signed(_T_375) & $signed(32'shf); // @[Math.scala 406:56:@33495.4]
  assign _T_378 = $signed(_T_377); // @[Math.scala 406:56:@33496.4]
  assign x420_sum_number = x420_sum_1_io_result; // @[Math.scala 154:22:@33507.4 Math.scala 155:14:@33508.4]
  assign _T_385 = x420_sum_number[31]; // @[FixedPoint.scala 50:25:@33512.4]
  assign _T_389 = _T_385 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33514.4]
  assign _T_390 = x420_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33515.4]
  assign _T_396 = _T_390 == 30'h3fffffff; // @[Math.scala 451:55:@33517.4]
  assign _T_397 = x420_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33518.4]
  assign _T_403 = _T_397 != 2'h0; // @[Math.scala 451:110:@33520.4]
  assign _T_404 = _T_396 & _T_403; // @[Math.scala 451:94:@33521.4]
  assign _T_406 = {_T_389,_T_390}; // @[Cat.scala 30:58:@33523.4]
  assign _T_416 = $signed(x420_sum_number); // @[Math.scala 406:49:@33531.4]
  assign _T_418 = $signed(_T_416) & $signed(32'sh3); // @[Math.scala 406:56:@33533.4]
  assign _T_419 = $signed(_T_418); // @[Math.scala 406:56:@33534.4]
  assign x423_sum_number = x423_sum_1_io_result; // @[Math.scala 154:22:@33545.4 Math.scala 155:14:@33546.4]
  assign _T_426 = x423_sum_number[31]; // @[FixedPoint.scala 50:25:@33550.4]
  assign _T_430 = _T_426 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33552.4]
  assign _T_431 = x423_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33553.4]
  assign _T_437 = _T_431 == 30'h3fffffff; // @[Math.scala 451:55:@33555.4]
  assign _T_438 = x423_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33556.4]
  assign _T_444 = _T_438 != 2'h0; // @[Math.scala 451:110:@33558.4]
  assign _T_445 = _T_437 & _T_444; // @[Math.scala 451:94:@33559.4]
  assign _T_449 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33567.4 package.scala 96:25:@33568.4]
  assign _T_459 = $signed(x423_sum_number); // @[Math.scala 406:49:@33576.4]
  assign _T_461 = $signed(_T_459) & $signed(32'sh3); // @[Math.scala 406:56:@33578.4]
  assign _T_462 = $signed(_T_461); // @[Math.scala 406:56:@33579.4]
  assign _T_466 = $signed(RetimeWrapper_2_io_out); // @[package.scala 96:25:@33587.4]
  assign x426_sum_number = x426_sum_1_io_result; // @[Math.scala 154:22:@33599.4 Math.scala 155:14:@33600.4]
  assign _T_473 = x426_sum_number[31]; // @[FixedPoint.scala 50:25:@33604.4]
  assign _T_477 = _T_473 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33606.4]
  assign _T_478 = x426_sum_number[31:2]; // @[FixedPoint.scala 18:52:@33607.4]
  assign _T_484 = _T_478 == 30'h3fffffff; // @[Math.scala 451:55:@33609.4]
  assign _T_485 = x426_sum_number[1:0]; // @[FixedPoint.scala 18:52:@33610.4]
  assign _T_491 = _T_485 != 2'h0; // @[Math.scala 451:110:@33612.4]
  assign _T_492 = _T_484 & _T_491; // @[Math.scala 451:94:@33613.4]
  assign _T_494 = {_T_477,_T_478}; // @[Cat.scala 30:58:@33615.4]
  assign _T_504 = $signed(x426_sum_number); // @[Math.scala 406:49:@33623.4]
  assign _T_506 = $signed(_T_504) & $signed(32'sh3); // @[Math.scala 406:56:@33625.4]
  assign _T_507 = $signed(_T_506); // @[Math.scala 406:56:@33626.4]
  assign x429_sum_number = x429_sum_1_io_result; // @[Math.scala 154:22:@33637.4 Math.scala 155:14:@33638.4]
  assign _T_517 = $signed(x429_sum_number); // @[Math.scala 476:37:@33643.4]
  assign x498_x430_D1 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@33681.4 package.scala 96:25:@33682.4]
  assign x499_x429_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@33690.4 package.scala 96:25:@33691.4]
  assign x432_sub_number = x432_sub_1_io_result; // @[Math.scala 195:22:@33663.4 Math.scala 196:14:@33664.4]
  assign _T_548 = x410_number[31]; // @[FixedPoint.scala 50:25:@33698.4]
  assign _T_552 = _T_548 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33700.4]
  assign _T_553 = x410_number[31:2]; // @[FixedPoint.scala 18:52:@33701.4]
  assign _T_559 = _T_553 == 30'h3fffffff; // @[Math.scala 451:55:@33703.4]
  assign _T_560 = x410_number[1:0]; // @[FixedPoint.scala 18:52:@33704.4]
  assign _T_566 = _T_560 != 2'h0; // @[Math.scala 451:110:@33706.4]
  assign _T_567 = _T_559 & _T_566; // @[Math.scala 451:94:@33707.4]
  assign _T_569 = {_T_552,_T_553}; // @[Cat.scala 30:58:@33709.4]
  assign x240_1_number = _T_567 ? 32'h0 : _T_569; // @[Math.scala 454:20:@33710.4]
  assign _GEN_0 = {{9'd0}, x240_1_number}; // @[Math.scala 461:32:@33715.4]
  assign _T_574 = _GEN_0 << 9; // @[Math.scala 461:32:@33715.4]
  assign _GEN_1 = {{7'd0}, x240_1_number}; // @[Math.scala 461:32:@33720.4]
  assign _T_577 = _GEN_1 << 7; // @[Math.scala 461:32:@33720.4]
  assign _T_610 = ~ io_sigsIn_break; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:101:@33809.4]
  assign _T_614 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@33817.4 package.scala 96:25:@33818.4]
  assign _T_616 = io_rr ? _T_614 : 1'h0; // @[implicits.scala 55:10:@33819.4]
  assign _T_617 = _T_610 & _T_616; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:118:@33820.4]
  assign _T_619 = _T_617 & _T_610; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:207:@33822.4]
  assign _T_620 = _T_619 & io_sigsIn_backpressure; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:226:@33823.4]
  assign x502_b229_D21 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@33779.4 package.scala 96:25:@33780.4]
  assign _T_621 = _T_620 & x502_b229_D21; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 164:252:@33824.4]
  assign x504_b230_D21 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@33797.4 package.scala 96:25:@33798.4]
  assign x506_b227_D23_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@33838.4 package.scala 96:25:@33839.4]
  assign _T_633 = $signed(x506_b227_D23_number); // @[Math.scala 476:37:@33846.4]
  assign x507_b228_D23_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@33863.4 package.scala 96:25:@33864.4]
  assign _T_646 = $signed(x507_b228_D23_number); // @[Math.scala 476:37:@33869.4]
  assign x246 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@33854.4 package.scala 96:25:@33855.4]
  assign x247 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@33877.4 package.scala 96:25:@33878.4]
  assign x248 = x246 | x247; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 183:24:@33881.4]
  assign _T_684 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@33949.4 package.scala 96:25:@33950.4]
  assign _T_686 = io_rr ? _T_684 : 1'h0; // @[implicits.scala 55:10:@33951.4]
  assign _T_687 = _T_610 & _T_686; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 202:194:@33952.4]
  assign x508_x249_D21 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@33892.4 package.scala 96:25:@33893.4]
  assign _T_688 = _T_687 & x508_x249_D21; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 202:283:@33953.4]
  assign x511_b229_D45 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@33919.4 package.scala 96:25:@33920.4]
  assign _T_689 = _T_688 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 202:291:@33954.4]
  assign x512_b230_D45 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@33928.4 package.scala 96:25:@33929.4]
  assign x252_rdcol_number = x252_rdcol_1_io_result; // @[Math.scala 195:22:@33973.4 Math.scala 196:14:@33974.4]
  assign _T_704 = $signed(x252_rdcol_number); // @[Math.scala 476:37:@33979.4]
  assign x514_x246_D1 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@33996.4 package.scala 96:25:@33997.4]
  assign x253 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@33987.4 package.scala 96:25:@33988.4]
  assign x254 = x514_x246_D1 | x253; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 212:24:@34000.4]
  assign _T_718 = x252_rdcol_number[31]; // @[FixedPoint.scala 50:25:@34007.4]
  assign _T_722 = _T_718 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@34009.4]
  assign _T_723 = x252_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@34010.4]
  assign _T_729 = _T_723 == 16'hffff; // @[Math.scala 451:55:@34012.4]
  assign _T_730 = x252_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@34013.4]
  assign _T_736 = _T_730 != 16'h0; // @[Math.scala 451:110:@34015.4]
  assign _T_737 = _T_729 & _T_736; // @[Math.scala 451:94:@34016.4]
  assign _T_739 = {_T_722,_T_723}; // @[Cat.scala 30:58:@34018.4]
  assign _T_751 = $signed(_T_704) & $signed(32'shffff); // @[Math.scala 406:56:@34028.4]
  assign _T_752 = $signed(_T_751); // @[Math.scala 406:56:@34029.4]
  assign x439_sum_number = x439_sum_1_io_result; // @[Math.scala 154:22:@34040.4 Math.scala 155:14:@34041.4]
  assign _T_759 = x439_sum_number[31]; // @[FixedPoint.scala 50:25:@34045.4]
  assign _T_763 = _T_759 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@34047.4]
  assign _T_764 = x439_sum_number[31:8]; // @[FixedPoint.scala 18:52:@34048.4]
  assign _T_770 = _T_764 == 24'hffffff; // @[Math.scala 451:55:@34050.4]
  assign _T_771 = x439_sum_number[7:0]; // @[FixedPoint.scala 18:52:@34051.4]
  assign _T_777 = _T_771 != 8'h0; // @[Math.scala 451:110:@34053.4]
  assign _T_778 = _T_770 & _T_777; // @[Math.scala 451:94:@34054.4]
  assign _T_782 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@34062.4 package.scala 96:25:@34063.4]
  assign _T_792 = $signed(x439_sum_number); // @[Math.scala 406:49:@34071.4]
  assign _T_794 = $signed(_T_792) & $signed(32'shff); // @[Math.scala 406:56:@34073.4]
  assign _T_795 = $signed(_T_794); // @[Math.scala 406:56:@34074.4]
  assign _T_799 = $signed(RetimeWrapper_27_io_out); // @[package.scala 96:25:@34082.4]
  assign x442_sum_number = x442_sum_1_io_result; // @[Math.scala 154:22:@34094.4 Math.scala 155:14:@34095.4]
  assign _T_806 = x442_sum_number[31]; // @[FixedPoint.scala 50:25:@34099.4]
  assign _T_810 = _T_806 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@34101.4]
  assign _T_811 = x442_sum_number[31:4]; // @[FixedPoint.scala 18:52:@34102.4]
  assign _T_817 = _T_811 == 28'hfffffff; // @[Math.scala 451:55:@34104.4]
  assign _T_818 = x442_sum_number[3:0]; // @[FixedPoint.scala 18:52:@34105.4]
  assign _T_824 = _T_818 != 4'h0; // @[Math.scala 451:110:@34107.4]
  assign _T_825 = _T_817 & _T_824; // @[Math.scala 451:94:@34108.4]
  assign _T_827 = {_T_810,_T_811}; // @[Cat.scala 30:58:@34110.4]
  assign _T_837 = $signed(x442_sum_number); // @[Math.scala 406:49:@34118.4]
  assign _T_839 = $signed(_T_837) & $signed(32'shf); // @[Math.scala 406:56:@34120.4]
  assign _T_840 = $signed(_T_839); // @[Math.scala 406:56:@34121.4]
  assign x445_sum_number = x445_sum_1_io_result; // @[Math.scala 154:22:@34132.4 Math.scala 155:14:@34133.4]
  assign _T_847 = x445_sum_number[31]; // @[FixedPoint.scala 50:25:@34137.4]
  assign _T_851 = _T_847 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34139.4]
  assign _T_852 = x445_sum_number[31:2]; // @[FixedPoint.scala 18:52:@34140.4]
  assign _T_858 = _T_852 == 30'h3fffffff; // @[Math.scala 451:55:@34142.4]
  assign _T_859 = x445_sum_number[1:0]; // @[FixedPoint.scala 18:52:@34143.4]
  assign _T_865 = _T_859 != 2'h0; // @[Math.scala 451:110:@34145.4]
  assign _T_866 = _T_858 & _T_865; // @[Math.scala 451:94:@34146.4]
  assign _T_868 = {_T_851,_T_852}; // @[Cat.scala 30:58:@34148.4]
  assign _T_878 = $signed(x445_sum_number); // @[Math.scala 406:49:@34156.4]
  assign _T_880 = $signed(_T_878) & $signed(32'sh3); // @[Math.scala 406:56:@34158.4]
  assign _T_881 = $signed(_T_880); // @[Math.scala 406:56:@34159.4]
  assign x448_sum_number = x448_sum_1_io_result; // @[Math.scala 154:22:@34170.4 Math.scala 155:14:@34171.4]
  assign _T_888 = x448_sum_number[31]; // @[FixedPoint.scala 50:25:@34175.4]
  assign _T_892 = _T_888 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34177.4]
  assign _T_893 = x448_sum_number[31:2]; // @[FixedPoint.scala 18:52:@34178.4]
  assign _T_899 = _T_893 == 30'h3fffffff; // @[Math.scala 451:55:@34180.4]
  assign _T_900 = x448_sum_number[1:0]; // @[FixedPoint.scala 18:52:@34181.4]
  assign _T_906 = _T_900 != 2'h0; // @[Math.scala 451:110:@34183.4]
  assign _T_907 = _T_899 & _T_906; // @[Math.scala 451:94:@34184.4]
  assign _T_909 = {_T_892,_T_893}; // @[Cat.scala 30:58:@34186.4]
  assign _T_919 = $signed(x448_sum_number); // @[Math.scala 406:49:@34194.4]
  assign _T_921 = $signed(_T_919) & $signed(32'sh3); // @[Math.scala 406:56:@34196.4]
  assign _T_922 = $signed(_T_921); // @[Math.scala 406:56:@34197.4]
  assign x451_sum_number = x451_sum_1_io_result; // @[Math.scala 154:22:@34208.4 Math.scala 155:14:@34209.4]
  assign _T_929 = x451_sum_number[31]; // @[FixedPoint.scala 50:25:@34213.4]
  assign _T_933 = _T_929 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34215.4]
  assign _T_934 = x451_sum_number[31:2]; // @[FixedPoint.scala 18:52:@34216.4]
  assign _T_940 = _T_934 == 30'h3fffffff; // @[Math.scala 451:55:@34218.4]
  assign _T_941 = x451_sum_number[1:0]; // @[FixedPoint.scala 18:52:@34219.4]
  assign _T_947 = _T_941 != 2'h0; // @[Math.scala 451:110:@34221.4]
  assign _T_948 = _T_940 & _T_947; // @[Math.scala 451:94:@34222.4]
  assign _T_950 = {_T_933,_T_934}; // @[Cat.scala 30:58:@34224.4]
  assign _T_960 = $signed(x451_sum_number); // @[Math.scala 406:49:@34232.4]
  assign _T_962 = $signed(_T_960) & $signed(32'sh3); // @[Math.scala 406:56:@34234.4]
  assign _T_963 = $signed(_T_962); // @[Math.scala 406:56:@34235.4]
  assign x454_sum_number = x454_sum_1_io_result; // @[Math.scala 154:22:@34246.4 Math.scala 155:14:@34247.4]
  assign _T_973 = $signed(x454_sum_number); // @[Math.scala 476:37:@34252.4]
  assign x455 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@34260.4 package.scala 96:25:@34261.4]
  assign x515_x454_sum_D1_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@34295.4 package.scala 96:25:@34296.4]
  assign x457_sub_number = x457_sub_1_io_result; // @[Math.scala 195:22:@34286.4 Math.scala 196:14:@34287.4]
  assign _T_1030 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@34359.4 package.scala 96:25:@34360.4]
  assign _T_1032 = io_rr ? _T_1030 : 1'h0; // @[implicits.scala 55:10:@34361.4]
  assign _T_1033 = _T_610 & _T_1032; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 275:194:@34362.4]
  assign x517_x255_D20 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@34338.4 package.scala 96:25:@34339.4]
  assign _T_1034 = _T_1033 & x517_x255_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 275:283:@34363.4]
  assign _T_1035 = _T_1034 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 275:291:@34364.4]
  assign x261_rdcol_number = x261_rdcol_1_io_result; // @[Math.scala 195:22:@34383.4 Math.scala 196:14:@34384.4]
  assign _T_1052 = $signed(x261_rdcol_number); // @[Math.scala 476:37:@34391.4]
  assign x262 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@34399.4 package.scala 96:25:@34400.4]
  assign x263 = x514_x246_D1 | x262; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 291:59:@34403.4]
  assign _T_1063 = x261_rdcol_number[31]; // @[FixedPoint.scala 50:25:@34410.4]
  assign _T_1067 = _T_1063 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@34412.4]
  assign _T_1068 = x261_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@34413.4]
  assign _T_1074 = _T_1068 == 16'hffff; // @[Math.scala 451:55:@34415.4]
  assign _T_1075 = x261_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@34416.4]
  assign _T_1081 = _T_1075 != 16'h0; // @[Math.scala 451:110:@34418.4]
  assign _T_1082 = _T_1074 & _T_1081; // @[Math.scala 451:94:@34419.4]
  assign _T_1084 = {_T_1067,_T_1068}; // @[Cat.scala 30:58:@34421.4]
  assign _T_1096 = $signed(_T_1052) & $signed(32'shffff); // @[Math.scala 406:56:@34431.4]
  assign _T_1097 = $signed(_T_1096); // @[Math.scala 406:56:@34432.4]
  assign x461_sum_number = x461_sum_1_io_result; // @[Math.scala 154:22:@34443.4 Math.scala 155:14:@34444.4]
  assign _T_1104 = x461_sum_number[31]; // @[FixedPoint.scala 50:25:@34448.4]
  assign _T_1108 = _T_1104 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@34450.4]
  assign _T_1109 = x461_sum_number[31:8]; // @[FixedPoint.scala 18:52:@34451.4]
  assign _T_1115 = _T_1109 == 24'hffffff; // @[Math.scala 451:55:@34453.4]
  assign _T_1116 = x461_sum_number[7:0]; // @[FixedPoint.scala 18:52:@34454.4]
  assign _T_1122 = _T_1116 != 8'h0; // @[Math.scala 451:110:@34456.4]
  assign _T_1123 = _T_1115 & _T_1122; // @[Math.scala 451:94:@34457.4]
  assign _T_1127 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@34465.4 package.scala 96:25:@34466.4]
  assign _T_1137 = $signed(x461_sum_number); // @[Math.scala 406:49:@34474.4]
  assign _T_1139 = $signed(_T_1137) & $signed(32'shff); // @[Math.scala 406:56:@34476.4]
  assign _T_1140 = $signed(_T_1139); // @[Math.scala 406:56:@34477.4]
  assign _T_1144 = $signed(RetimeWrapper_37_io_out); // @[package.scala 96:25:@34485.4]
  assign x464_sum_number = x464_sum_1_io_result; // @[Math.scala 154:22:@34497.4 Math.scala 155:14:@34498.4]
  assign _T_1151 = x464_sum_number[31]; // @[FixedPoint.scala 50:25:@34502.4]
  assign _T_1155 = _T_1151 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@34504.4]
  assign _T_1156 = x464_sum_number[31:4]; // @[FixedPoint.scala 18:52:@34505.4]
  assign _T_1162 = _T_1156 == 28'hfffffff; // @[Math.scala 451:55:@34507.4]
  assign _T_1163 = x464_sum_number[3:0]; // @[FixedPoint.scala 18:52:@34508.4]
  assign _T_1169 = _T_1163 != 4'h0; // @[Math.scala 451:110:@34510.4]
  assign _T_1170 = _T_1162 & _T_1169; // @[Math.scala 451:94:@34511.4]
  assign _T_1172 = {_T_1155,_T_1156}; // @[Cat.scala 30:58:@34513.4]
  assign _T_1182 = $signed(x464_sum_number); // @[Math.scala 406:49:@34521.4]
  assign _T_1184 = $signed(_T_1182) & $signed(32'shf); // @[Math.scala 406:56:@34523.4]
  assign _T_1185 = $signed(_T_1184); // @[Math.scala 406:56:@34524.4]
  assign x467_sum_number = x467_sum_1_io_result; // @[Math.scala 154:22:@34535.4 Math.scala 155:14:@34536.4]
  assign _T_1192 = x467_sum_number[31]; // @[FixedPoint.scala 50:25:@34540.4]
  assign _T_1196 = _T_1192 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34542.4]
  assign _T_1197 = x467_sum_number[31:2]; // @[FixedPoint.scala 18:52:@34543.4]
  assign _T_1203 = _T_1197 == 30'h3fffffff; // @[Math.scala 451:55:@34545.4]
  assign _T_1204 = x467_sum_number[1:0]; // @[FixedPoint.scala 18:52:@34546.4]
  assign _T_1210 = _T_1204 != 2'h0; // @[Math.scala 451:110:@34548.4]
  assign _T_1211 = _T_1203 & _T_1210; // @[Math.scala 451:94:@34549.4]
  assign _T_1213 = {_T_1196,_T_1197}; // @[Cat.scala 30:58:@34551.4]
  assign _T_1223 = $signed(x467_sum_number); // @[Math.scala 406:49:@34559.4]
  assign _T_1225 = $signed(_T_1223) & $signed(32'sh3); // @[Math.scala 406:56:@34561.4]
  assign _T_1226 = $signed(_T_1225); // @[Math.scala 406:56:@34562.4]
  assign x470_sum_number = x470_sum_1_io_result; // @[Math.scala 154:22:@34573.4 Math.scala 155:14:@34574.4]
  assign _T_1233 = x470_sum_number[31]; // @[FixedPoint.scala 50:25:@34578.4]
  assign _T_1237 = _T_1233 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34580.4]
  assign _T_1238 = x470_sum_number[31:2]; // @[FixedPoint.scala 18:52:@34581.4]
  assign _T_1244 = _T_1238 == 30'h3fffffff; // @[Math.scala 451:55:@34583.4]
  assign _T_1245 = x470_sum_number[1:0]; // @[FixedPoint.scala 18:52:@34584.4]
  assign _T_1251 = _T_1245 != 2'h0; // @[Math.scala 451:110:@34586.4]
  assign _T_1252 = _T_1244 & _T_1251; // @[Math.scala 451:94:@34587.4]
  assign _T_1254 = {_T_1237,_T_1238}; // @[Cat.scala 30:58:@34589.4]
  assign _T_1264 = $signed(x470_sum_number); // @[Math.scala 406:49:@34597.4]
  assign _T_1266 = $signed(_T_1264) & $signed(32'sh3); // @[Math.scala 406:56:@34599.4]
  assign _T_1267 = $signed(_T_1266); // @[Math.scala 406:56:@34600.4]
  assign x473_sum_number = x473_sum_1_io_result; // @[Math.scala 154:22:@34611.4 Math.scala 155:14:@34612.4]
  assign _T_1274 = x473_sum_number[31]; // @[FixedPoint.scala 50:25:@34616.4]
  assign _T_1278 = _T_1274 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34618.4]
  assign _T_1279 = x473_sum_number[31:2]; // @[FixedPoint.scala 18:52:@34619.4]
  assign _T_1285 = _T_1279 == 30'h3fffffff; // @[Math.scala 451:55:@34621.4]
  assign _T_1286 = x473_sum_number[1:0]; // @[FixedPoint.scala 18:52:@34622.4]
  assign _T_1292 = _T_1286 != 2'h0; // @[Math.scala 451:110:@34624.4]
  assign _T_1293 = _T_1285 & _T_1292; // @[Math.scala 451:94:@34625.4]
  assign _T_1295 = {_T_1278,_T_1279}; // @[Cat.scala 30:58:@34627.4]
  assign _T_1305 = $signed(x473_sum_number); // @[Math.scala 406:49:@34635.4]
  assign _T_1307 = $signed(_T_1305) & $signed(32'sh3); // @[Math.scala 406:56:@34637.4]
  assign _T_1308 = $signed(_T_1307); // @[Math.scala 406:56:@34638.4]
  assign x476_sum_number = x476_sum_1_io_result; // @[Math.scala 154:22:@34649.4 Math.scala 155:14:@34650.4]
  assign _T_1318 = $signed(x476_sum_number); // @[Math.scala 476:37:@34655.4]
  assign x477 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@34663.4 package.scala 96:25:@34664.4]
  assign x519_x476_sum_D1_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@34698.4 package.scala 96:25:@34699.4]
  assign x479_sub_number = x479_sub_1_io_result; // @[Math.scala 195:22:@34689.4 Math.scala 196:14:@34690.4]
  assign _T_1372 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@34753.4 package.scala 96:25:@34754.4]
  assign _T_1374 = io_rr ? _T_1372 : 1'h0; // @[implicits.scala 55:10:@34755.4]
  assign _T_1375 = _T_610 & _T_1374; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 352:194:@34756.4]
  assign x521_x264_D20 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@34741.4 package.scala 96:25:@34742.4]
  assign _T_1376 = _T_1375 & x521_x264_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 352:283:@34757.4]
  assign _T_1377 = _T_1376 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 352:291:@34758.4]
  assign x270_rdrow_number = x270_rdrow_1_io_result; // @[Math.scala 195:22:@34777.4 Math.scala 196:14:@34778.4]
  assign _T_1394 = $signed(x270_rdrow_number); // @[Math.scala 406:49:@34784.4]
  assign _T_1396 = $signed(_T_1394) & $signed(32'sh3); // @[Math.scala 406:56:@34786.4]
  assign _T_1397 = $signed(_T_1396); // @[Math.scala 406:56:@34787.4]
  assign x481_number = $unsigned(_T_1397); // @[implicits.scala 133:21:@34788.4]
  assign x272 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@34802.4 package.scala 96:25:@34803.4]
  assign x522_x247_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@34811.4 package.scala 96:25:@34812.4]
  assign x273 = x272 | x522_x247_D1; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 364:24:@34815.4]
  assign _T_1423 = $signed(x481_number); // @[Math.scala 406:49:@34824.4]
  assign _T_1425 = $signed(_T_1423) & $signed(32'sh3); // @[Math.scala 406:56:@34826.4]
  assign _T_1426 = $signed(_T_1425); // @[Math.scala 406:56:@34827.4]
  assign _T_1430 = $signed(RetimeWrapper_46_io_out); // @[package.scala 96:25:@34835.4]
  assign _T_1434 = x481_number[31]; // @[FixedPoint.scala 50:25:@34842.4]
  assign _T_1438 = _T_1434 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34844.4]
  assign _T_1439 = x481_number[31:2]; // @[FixedPoint.scala 18:52:@34845.4]
  assign _T_1445 = _T_1439 == 30'h3fffffff; // @[Math.scala 451:55:@34847.4]
  assign _T_1446 = x481_number[1:0]; // @[FixedPoint.scala 18:52:@34848.4]
  assign _T_1452 = _T_1446 != 2'h0; // @[Math.scala 451:110:@34850.4]
  assign _T_1453 = _T_1445 & _T_1452; // @[Math.scala 451:94:@34851.4]
  assign _T_1457 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@34859.4 package.scala 96:25:@34860.4]
  assign x276_1_number = _T_1453 ? 32'h0 : _T_1457; // @[Math.scala 454:20:@34861.4]
  assign _GEN_2 = {{9'd0}, x276_1_number}; // @[Math.scala 461:32:@34866.4]
  assign _T_1462 = _GEN_2 << 9; // @[Math.scala 461:32:@34866.4]
  assign _GEN_3 = {{7'd0}, x276_1_number}; // @[Math.scala 461:32:@34871.4]
  assign _T_1465 = _GEN_3 << 7; // @[Math.scala 461:32:@34871.4]
  assign _T_1498 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@34948.4 package.scala 96:25:@34949.4]
  assign _T_1500 = io_rr ? _T_1498 : 1'h0; // @[implicits.scala 55:10:@34950.4]
  assign _T_1501 = _T_610 & _T_1500; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 399:194:@34951.4]
  assign x525_x274_D20 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@34918.4 package.scala 96:25:@34919.4]
  assign _T_1502 = _T_1501 & x525_x274_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 399:283:@34952.4]
  assign _T_1503 = _T_1502 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 399:326:@34953.4]
  assign x281 = x272 | x253; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 403:59:@34964.4]
  assign _T_1532 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@35008.4 package.scala 96:25:@35009.4]
  assign _T_1534 = io_rr ? _T_1532 : 1'h0; // @[implicits.scala 55:10:@35010.4]
  assign _T_1535 = _T_610 & _T_1534; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 418:194:@35011.4]
  assign x529_x282_D20 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@34996.4 package.scala 96:25:@34997.4]
  assign _T_1536 = _T_1535 & x529_x282_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 418:283:@35012.4]
  assign _T_1537 = _T_1536 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 418:291:@35013.4]
  assign x286 = x272 | x262; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 422:59:@35024.4]
  assign _T_1561 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@35057.4 package.scala 96:25:@35058.4]
  assign _T_1563 = io_rr ? _T_1561 : 1'h0; // @[implicits.scala 55:10:@35059.4]
  assign _T_1564 = _T_610 & _T_1563; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 433:194:@35060.4]
  assign x530_x287_D20 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@35045.4 package.scala 96:25:@35046.4]
  assign _T_1565 = _T_1564 & x530_x287_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 433:283:@35061.4]
  assign _T_1566 = _T_1565 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 433:291:@35062.4]
  assign x291_rdrow_number = x291_rdrow_1_io_result; // @[Math.scala 195:22:@35081.4 Math.scala 196:14:@35082.4]
  assign _T_1583 = $signed(x291_rdrow_number); // @[Math.scala 406:49:@35088.4]
  assign _T_1585 = $signed(_T_1583) & $signed(32'sh3); // @[Math.scala 406:56:@35090.4]
  assign _T_1586 = $signed(_T_1585); // @[Math.scala 406:56:@35091.4]
  assign x486_number = $unsigned(_T_1586); // @[implicits.scala 133:21:@35092.4]
  assign x293 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@35106.4 package.scala 96:25:@35107.4]
  assign x294 = x293 | x522_x247_D1; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 443:24:@35110.4]
  assign _T_1609 = $signed(x486_number); // @[Math.scala 406:49:@35119.4]
  assign _T_1611 = $signed(_T_1609) & $signed(32'sh3); // @[Math.scala 406:56:@35121.4]
  assign _T_1612 = $signed(_T_1611); // @[Math.scala 406:56:@35122.4]
  assign _T_1616 = $signed(RetimeWrapper_60_io_out); // @[package.scala 96:25:@35130.4]
  assign _T_1620 = x486_number[31]; // @[FixedPoint.scala 50:25:@35137.4]
  assign _T_1624 = _T_1620 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@35139.4]
  assign _T_1625 = x486_number[31:2]; // @[FixedPoint.scala 18:52:@35140.4]
  assign _T_1631 = _T_1625 == 30'h3fffffff; // @[Math.scala 451:55:@35142.4]
  assign _T_1632 = x486_number[1:0]; // @[FixedPoint.scala 18:52:@35143.4]
  assign _T_1638 = _T_1632 != 2'h0; // @[Math.scala 451:110:@35145.4]
  assign _T_1639 = _T_1631 & _T_1638; // @[Math.scala 451:94:@35146.4]
  assign _T_1643 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@35154.4 package.scala 96:25:@35155.4]
  assign x297_1_number = _T_1639 ? 32'h0 : _T_1643; // @[Math.scala 454:20:@35156.4]
  assign _GEN_4 = {{9'd0}, x297_1_number}; // @[Math.scala 461:32:@35161.4]
  assign _T_1648 = _GEN_4 << 9; // @[Math.scala 461:32:@35161.4]
  assign _GEN_5 = {{7'd0}, x297_1_number}; // @[Math.scala 461:32:@35166.4]
  assign _T_1651 = _GEN_5 << 7; // @[Math.scala 461:32:@35166.4]
  assign _T_1681 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@35234.4 package.scala 96:25:@35235.4]
  assign _T_1683 = io_rr ? _T_1681 : 1'h0; // @[implicits.scala 55:10:@35236.4]
  assign _T_1684 = _T_610 & _T_1683; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 470:194:@35237.4]
  assign x534_x295_D20 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@35222.4 package.scala 96:25:@35223.4]
  assign _T_1685 = _T_1684 & x534_x295_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 470:283:@35238.4]
  assign _T_1686 = _T_1685 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 470:291:@35239.4]
  assign x302 = x293 | x253; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 474:24:@35250.4]
  assign _T_1713 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@35292.4 package.scala 96:25:@35293.4]
  assign _T_1715 = io_rr ? _T_1713 : 1'h0; // @[implicits.scala 55:10:@35294.4]
  assign _T_1716 = _T_610 & _T_1715; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 487:194:@35295.4]
  assign x536_x303_D20 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@35280.4 package.scala 96:25:@35281.4]
  assign _T_1717 = _T_1716 & x536_x303_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 487:283:@35296.4]
  assign _T_1718 = _T_1717 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 487:291:@35297.4]
  assign x307 = x293 | x262; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 491:24:@35308.4]
  assign _T_1742 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@35341.4 package.scala 96:25:@35342.4]
  assign _T_1744 = io_rr ? _T_1742 : 1'h0; // @[implicits.scala 55:10:@35343.4]
  assign _T_1745 = _T_610 & _T_1744; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 502:194:@35344.4]
  assign x537_x308_D20 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@35329.4 package.scala 96:25:@35330.4]
  assign _T_1746 = _T_1745 & x537_x308_D20; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 502:283:@35345.4]
  assign _T_1747 = _T_1746 & x511_b229_D45; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 502:291:@35346.4]
  assign _T_1878 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@35647.4 package.scala 96:25:@35648.4]
  assign _T_1880 = io_rr ? _T_1878 : 1'h0; // @[implicits.scala 55:10:@35649.4]
  assign _T_1881 = _T_610 & _T_1880; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:167:@35650.4]
  assign _T_1883 = _T_1881 & _T_610; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:256:@35652.4]
  assign _T_1884 = _T_1883 & io_sigsIn_backpressure; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:275:@35653.4]
  assign x541_b229_D64 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@35609.4 package.scala 96:25:@35610.4]
  assign _T_1885 = _T_1884 & x541_b229_D64; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 572:301:@35654.4]
  assign x542_b230_D64 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@35618.4 package.scala 96:25:@35619.4]
  assign _T_1916 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@35725.4 package.scala 96:25:@35726.4]
  assign _T_1918 = io_rr ? _T_1916 : 1'h0; // @[implicits.scala 55:10:@35727.4]
  assign _T_1919 = _T_610 & _T_1918; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 590:195:@35728.4]
  assign x545_x249_D41 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@35668.4 package.scala 96:25:@35669.4]
  assign _T_1920 = _T_1919 & x545_x249_D41; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 590:284:@35729.4]
  assign x548_b229_D65 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@35695.4 package.scala 96:25:@35696.4]
  assign _T_1921 = _T_1920 & x548_b229_D65; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 590:292:@35730.4]
  assign x549_b230_D65 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@35704.4 package.scala 96:25:@35705.4]
  assign _T_1944 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@35776.4 package.scala 96:25:@35777.4]
  assign _T_1946 = io_rr ? _T_1944 : 1'h0; // @[implicits.scala 55:10:@35778.4]
  assign _T_1947 = _T_610 & _T_1946; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 603:195:@35779.4]
  assign x551_x255_D40 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@35746.4 package.scala 96:25:@35747.4]
  assign _T_1948 = _T_1947 & x551_x255_D40; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 603:284:@35780.4]
  assign _T_1949 = _T_1948 & x548_b229_D65; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 603:292:@35781.4]
  assign _T_1972 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@35827.4 package.scala 96:25:@35828.4]
  assign _T_1974 = io_rr ? _T_1972 : 1'h0; // @[implicits.scala 55:10:@35829.4]
  assign _T_1975 = _T_610 & _T_1974; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 616:195:@35830.4]
  assign x554_x274_D40 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@35797.4 package.scala 96:25:@35798.4]
  assign _T_1976 = _T_1975 & x554_x274_D40; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 616:284:@35831.4]
  assign _T_1977 = _T_1976 & x548_b229_D65; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 616:292:@35832.4]
  assign _T_1997 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@35869.4 package.scala 96:25:@35870.4]
  assign _T_1999 = io_rr ? _T_1997 : 1'h0; // @[implicits.scala 55:10:@35871.4]
  assign _T_2000 = _T_610 & _T_1999; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 627:195:@35872.4]
  assign x557_x282_D40 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@35848.4 package.scala 96:25:@35849.4]
  assign _T_2001 = _T_2000 & x557_x282_D40; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 627:284:@35873.4]
  assign _T_2002 = _T_2001 & x548_b229_D65; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 627:292:@35874.4]
  assign _T_2076 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@36031.4 package.scala 96:25:@36032.4]
  assign _T_2078 = io_rr ? _T_2076 : 1'h0; // @[implicits.scala 55:10:@36033.4]
  assign x560_b229_D84 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@36022.4 package.scala 96:25:@36023.4]
  assign _T_2079 = _T_2078 & x560_b229_D84; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 667:117:@36034.4]
  assign x559_b230_D84 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@36013.4 package.scala 96:25:@36014.4]
  assign _T_2080 = _T_2079 & x559_b230_D84; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 667:123:@36035.4]
  assign x243_sum_number = x243_sum_1_io_result; // @[Math.scala 154:22:@33761.4 Math.scala 155:14:@33762.4]
  assign x501_x411_D21_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@33770.4 package.scala 96:25:@33771.4]
  assign x505_x433_D13_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@33806.4 package.scala 96:25:@33807.4]
  assign x509_x411_D45_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@33901.4 package.scala 96:25:@33902.4]
  assign x510_x243_sum_D24_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@33910.4 package.scala 96:25:@33911.4]
  assign x513_x433_D37_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@33937.4 package.scala 96:25:@33938.4]
  assign x258_sum_number = x258_sum_1_io_result; // @[Math.scala 154:22:@34329.4 Math.scala 155:14:@34330.4]
  assign x518_x458_D13_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@34347.4 package.scala 96:25:@34348.4]
  assign x267_sum_number = x267_sum_1_io_result; // @[Math.scala 154:22:@34723.4 Math.scala 155:14:@34724.4]
  assign x520_x480_D13_number = RetimeWrapper_41_io_out; // @[package.scala 96:25:@34732.4 package.scala 96:25:@34733.4]
  assign x526_x278_sum_D1_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@34927.4 package.scala 96:25:@34928.4]
  assign x527_x482_D20_number = RetimeWrapper_52_io_out; // @[package.scala 96:25:@34936.4 package.scala 96:25:@34937.4]
  assign x283_sum_number = x283_sum_1_io_result; // @[Math.scala 154:22:@34987.4 Math.scala 155:14:@34988.4]
  assign x288_sum_number = x288_sum_1_io_result; // @[Math.scala 154:22:@35036.4 Math.scala 155:14:@35037.4]
  assign x532_x299_sum_D1_number = RetimeWrapper_63_io_out; // @[package.scala 96:25:@35204.4 package.scala 96:25:@35205.4]
  assign x533_x487_D20_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@35213.4 package.scala 96:25:@35214.4]
  assign x304_sum_number = x304_sum_1_io_result; // @[Math.scala 154:22:@35271.4 Math.scala 155:14:@35272.4]
  assign x309_sum_number = x309_sum_1_io_result; // @[Math.scala 154:22:@35320.4 Math.scala 155:14:@35321.4]
  assign x539_x411_D64_number = RetimeWrapper_73_io_out; // @[package.scala 96:25:@35591.4 package.scala 96:25:@35592.4]
  assign x540_x243_sum_D43_number = RetimeWrapper_74_io_out; // @[package.scala 96:25:@35600.4 package.scala 96:25:@35601.4]
  assign x544_x433_D56_number = RetimeWrapper_78_io_out; // @[package.scala 96:25:@35636.4 package.scala 96:25:@35637.4]
  assign x546_x411_D65_number = RetimeWrapper_81_io_out; // @[package.scala 96:25:@35677.4 package.scala 96:25:@35678.4]
  assign x547_x243_sum_D44_number = RetimeWrapper_82_io_out; // @[package.scala 96:25:@35686.4 package.scala 96:25:@35687.4]
  assign x550_x433_D57_number = RetimeWrapper_85_io_out; // @[package.scala 96:25:@35713.4 package.scala 96:25:@35714.4]
  assign x552_x458_D33_number = RetimeWrapper_88_io_out; // @[package.scala 96:25:@35755.4 package.scala 96:25:@35756.4]
  assign x553_x258_sum_D20_number = RetimeWrapper_89_io_out; // @[package.scala 96:25:@35764.4 package.scala 96:25:@35765.4]
  assign x555_x278_sum_D21_number = RetimeWrapper_92_io_out; // @[package.scala 96:25:@35806.4 package.scala 96:25:@35807.4]
  assign x556_x482_D40_number = RetimeWrapper_93_io_out; // @[package.scala 96:25:@35815.4 package.scala 96:25:@35816.4]
  assign x558_x283_sum_D20_number = RetimeWrapper_96_io_out; // @[package.scala 96:25:@35857.4 package.scala 96:25:@35858.4]
  assign io_in_x202_TVALID = _T_2080 & io_sigsIn_backpressure; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 667:22:@36037.4]
  assign io_in_x202_TDATA = {{224'd0}, RetimeWrapper_98_io_out}; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 668:24:@36038.4]
  assign io_in_x201_TREADY = _T_211 & _T_213; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 67:22:@33243.4 sm_x357_inr_Foreach_SAMPLER_BOX.scala 69:22:@33251.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@33221.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@33233.4]
  assign RetimeWrapper_clock = clock; // @[:@33254.4]
  assign RetimeWrapper_reset = reset; // @[:@33255.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33257.4]
  assign RetimeWrapper_io_in = io_in_x201_TDATA[31:0]; // @[package.scala 94:16:@33256.4]
  assign x233_lb_0_clock = clock; // @[:@33264.4]
  assign x233_lb_0_reset = reset; // @[:@33265.4]
  assign x233_lb_0_io_rPort_8_banks_1 = x520_x480_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@34761.4]
  assign x233_lb_0_io_rPort_8_banks_0 = x509_x411_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@34760.4]
  assign x233_lb_0_io_rPort_8_ofs_0 = x267_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@34762.4]
  assign x233_lb_0_io_rPort_8_en_0 = _T_1377 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@34764.4]
  assign x233_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34763.4]
  assign x233_lb_0_io_rPort_7_banks_1 = x518_x458_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@35300.4]
  assign x233_lb_0_io_rPort_7_banks_0 = x533_x487_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@35299.4]
  assign x233_lb_0_io_rPort_7_ofs_0 = x304_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@35301.4]
  assign x233_lb_0_io_rPort_7_en_0 = _T_1718 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@35303.4]
  assign x233_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35302.4]
  assign x233_lb_0_io_rPort_6_banks_1 = x513_x433_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@35242.4]
  assign x233_lb_0_io_rPort_6_banks_0 = x533_x487_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@35241.4]
  assign x233_lb_0_io_rPort_6_ofs_0 = x532_x299_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@35243.4]
  assign x233_lb_0_io_rPort_6_en_0 = _T_1686 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@35245.4]
  assign x233_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35244.4]
  assign x233_lb_0_io_rPort_5_banks_1 = x513_x433_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@33957.4]
  assign x233_lb_0_io_rPort_5_banks_0 = x509_x411_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@33956.4]
  assign x233_lb_0_io_rPort_5_ofs_0 = x510_x243_sum_D24_number[9:0]; // @[MemInterfaceType.scala 107:54:@33958.4]
  assign x233_lb_0_io_rPort_5_en_0 = _T_689 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@33960.4]
  assign x233_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33959.4]
  assign x233_lb_0_io_rPort_4_banks_1 = x520_x480_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@35349.4]
  assign x233_lb_0_io_rPort_4_banks_0 = x533_x487_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@35348.4]
  assign x233_lb_0_io_rPort_4_ofs_0 = x309_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@35350.4]
  assign x233_lb_0_io_rPort_4_en_0 = _T_1747 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@35352.4]
  assign x233_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35351.4]
  assign x233_lb_0_io_rPort_3_banks_1 = x518_x458_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@34367.4]
  assign x233_lb_0_io_rPort_3_banks_0 = x509_x411_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@34366.4]
  assign x233_lb_0_io_rPort_3_ofs_0 = x258_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@34368.4]
  assign x233_lb_0_io_rPort_3_en_0 = _T_1035 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@34370.4]
  assign x233_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34369.4]
  assign x233_lb_0_io_rPort_2_banks_1 = x513_x433_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@34956.4]
  assign x233_lb_0_io_rPort_2_banks_0 = x527_x482_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@34955.4]
  assign x233_lb_0_io_rPort_2_ofs_0 = x526_x278_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@34957.4]
  assign x233_lb_0_io_rPort_2_en_0 = _T_1503 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@34959.4]
  assign x233_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34958.4]
  assign x233_lb_0_io_rPort_1_banks_1 = x520_x480_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@35065.4]
  assign x233_lb_0_io_rPort_1_banks_0 = x527_x482_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@35064.4]
  assign x233_lb_0_io_rPort_1_ofs_0 = x288_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@35066.4]
  assign x233_lb_0_io_rPort_1_en_0 = _T_1566 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@35068.4]
  assign x233_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35067.4]
  assign x233_lb_0_io_rPort_0_banks_1 = x518_x458_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@35016.4]
  assign x233_lb_0_io_rPort_0_banks_0 = x527_x482_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@35015.4]
  assign x233_lb_0_io_rPort_0_ofs_0 = x283_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@35017.4]
  assign x233_lb_0_io_rPort_0_en_0 = _T_1537 & x512_b230_D45; // @[MemInterfaceType.scala 110:79:@35019.4]
  assign x233_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35018.4]
  assign x233_lb_0_io_wPort_0_banks_1 = x505_x433_D13_number[1:0]; // @[MemInterfaceType.scala 88:58:@33827.4]
  assign x233_lb_0_io_wPort_0_banks_0 = x501_x411_D21_number[2:0]; // @[MemInterfaceType.scala 88:58:@33826.4]
  assign x233_lb_0_io_wPort_0_ofs_0 = x243_sum_number[9:0]; // @[MemInterfaceType.scala 89:54:@33828.4]
  assign x233_lb_0_io_wPort_0_data_0 = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 90:56:@33829.4]
  assign x233_lb_0_io_wPort_0_en_0 = _T_621 & x504_b230_D21; // @[MemInterfaceType.scala 93:57:@33831.4]
  assign x234_lb2_0_clock = clock; // @[:@33331.4]
  assign x234_lb2_0_reset = reset; // @[:@33332.4]
  assign x234_lb2_0_io_rPort_3_banks_1 = x552_x458_D33_number[1:0]; // @[MemInterfaceType.scala 106:58:@35877.4]
  assign x234_lb2_0_io_rPort_3_banks_0 = x556_x482_D40_number[2:0]; // @[MemInterfaceType.scala 106:58:@35876.4]
  assign x234_lb2_0_io_rPort_3_ofs_0 = x558_x283_sum_D20_number[9:0]; // @[MemInterfaceType.scala 107:54:@35878.4]
  assign x234_lb2_0_io_rPort_3_en_0 = _T_2002 & x549_b230_D65; // @[MemInterfaceType.scala 110:79:@35880.4]
  assign x234_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35879.4]
  assign x234_lb2_0_io_rPort_2_banks_1 = x550_x433_D57_number[1:0]; // @[MemInterfaceType.scala 106:58:@35835.4]
  assign x234_lb2_0_io_rPort_2_banks_0 = x556_x482_D40_number[2:0]; // @[MemInterfaceType.scala 106:58:@35834.4]
  assign x234_lb2_0_io_rPort_2_ofs_0 = x555_x278_sum_D21_number[9:0]; // @[MemInterfaceType.scala 107:54:@35836.4]
  assign x234_lb2_0_io_rPort_2_en_0 = _T_1977 & x549_b230_D65; // @[MemInterfaceType.scala 110:79:@35838.4]
  assign x234_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35837.4]
  assign x234_lb2_0_io_rPort_1_banks_1 = x552_x458_D33_number[1:0]; // @[MemInterfaceType.scala 106:58:@35784.4]
  assign x234_lb2_0_io_rPort_1_banks_0 = x546_x411_D65_number[2:0]; // @[MemInterfaceType.scala 106:58:@35783.4]
  assign x234_lb2_0_io_rPort_1_ofs_0 = x553_x258_sum_D20_number[9:0]; // @[MemInterfaceType.scala 107:54:@35785.4]
  assign x234_lb2_0_io_rPort_1_en_0 = _T_1949 & x549_b230_D65; // @[MemInterfaceType.scala 110:79:@35787.4]
  assign x234_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35786.4]
  assign x234_lb2_0_io_rPort_0_banks_1 = x550_x433_D57_number[1:0]; // @[MemInterfaceType.scala 106:58:@35733.4]
  assign x234_lb2_0_io_rPort_0_banks_0 = x546_x411_D65_number[2:0]; // @[MemInterfaceType.scala 106:58:@35732.4]
  assign x234_lb2_0_io_rPort_0_ofs_0 = x547_x243_sum_D44_number[9:0]; // @[MemInterfaceType.scala 107:54:@35734.4]
  assign x234_lb2_0_io_rPort_0_en_0 = _T_1921 & x549_b230_D65; // @[MemInterfaceType.scala 110:79:@35736.4]
  assign x234_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35735.4]
  assign x234_lb2_0_io_wPort_0_banks_1 = x544_x433_D56_number[1:0]; // @[MemInterfaceType.scala 88:58:@35657.4]
  assign x234_lb2_0_io_wPort_0_banks_0 = x539_x411_D64_number[2:0]; // @[MemInterfaceType.scala 88:58:@35656.4]
  assign x234_lb2_0_io_wPort_0_ofs_0 = x540_x243_sum_D43_number[9:0]; // @[MemInterfaceType.scala 89:54:@35658.4]
  assign x234_lb2_0_io_wPort_0_data_0 = RetimeWrapper_77_io_out; // @[MemInterfaceType.scala 90:56:@35659.4]
  assign x234_lb2_0_io_wPort_0_en_0 = _T_1885 & x542_b230_D64; // @[MemInterfaceType.scala 93:57:@35661.4]
  assign x414_sum_1_clock = clock; // @[:@33426.4]
  assign x414_sum_1_reset = reset; // @[:@33427.4]
  assign x414_sum_1_io_a = _T_281 ? 32'h0 : _T_283; // @[Math.scala 151:17:@33428.4]
  assign x414_sum_1_io_b = $unsigned(_T_296); // @[Math.scala 152:17:@33429.4]
  assign x414_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33430.4]
  assign x417_sum_1_clock = clock; // @[:@33464.4]
  assign x417_sum_1_reset = reset; // @[:@33465.4]
  assign x417_sum_1_io_a = _T_322 ? 32'h0 : _T_324; // @[Math.scala 151:17:@33466.4]
  assign x417_sum_1_io_b = $unsigned(_T_337); // @[Math.scala 152:17:@33467.4]
  assign x417_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33468.4]
  assign x420_sum_1_clock = clock; // @[:@33502.4]
  assign x420_sum_1_reset = reset; // @[:@33503.4]
  assign x420_sum_1_io_a = _T_363 ? 32'h0 : _T_365; // @[Math.scala 151:17:@33504.4]
  assign x420_sum_1_io_b = $unsigned(_T_378); // @[Math.scala 152:17:@33505.4]
  assign x420_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33506.4]
  assign x423_sum_1_clock = clock; // @[:@33540.4]
  assign x423_sum_1_reset = reset; // @[:@33541.4]
  assign x423_sum_1_io_a = _T_404 ? 32'h0 : _T_406; // @[Math.scala 151:17:@33542.4]
  assign x423_sum_1_io_b = $unsigned(_T_419); // @[Math.scala 152:17:@33543.4]
  assign x423_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33544.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33563.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33564.4]
  assign RetimeWrapper_1_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@33566.4]
  assign RetimeWrapper_1_io_in = {_T_430,_T_431}; // @[package.scala 94:16:@33565.4]
  assign RetimeWrapper_2_clock = clock; // @[:@33581.4]
  assign RetimeWrapper_2_reset = reset; // @[:@33582.4]
  assign RetimeWrapper_2_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@33585.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_462); // @[package.scala 94:16:@33584.4]
  assign x426_sum_1_clock = clock; // @[:@33594.4]
  assign x426_sum_1_reset = reset; // @[:@33595.4]
  assign x426_sum_1_io_a = _T_445 ? 32'h0 : _T_449; // @[Math.scala 151:17:@33596.4]
  assign x426_sum_1_io_b = $unsigned(_T_466); // @[Math.scala 152:17:@33597.4]
  assign x426_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33598.4]
  assign x429_sum_1_clock = clock; // @[:@33632.4]
  assign x429_sum_1_reset = reset; // @[:@33633.4]
  assign x429_sum_1_io_a = _T_492 ? 32'h0 : _T_494; // @[Math.scala 151:17:@33634.4]
  assign x429_sum_1_io_b = $unsigned(_T_507); // @[Math.scala 152:17:@33635.4]
  assign x429_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33636.4]
  assign x432_sub_1_clock = clock; // @[:@33658.4]
  assign x432_sub_1_reset = reset; // @[:@33659.4]
  assign x432_sub_1_io_a = x429_sum_1_io_result; // @[Math.scala 192:17:@33660.4]
  assign x432_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@33661.4]
  assign x432_sub_1_io_flow = io_in_x202_TREADY; // @[Math.scala 194:20:@33662.4]
  assign RetimeWrapper_3_clock = clock; // @[:@33668.4]
  assign RetimeWrapper_3_reset = reset; // @[:@33669.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33671.4]
  assign RetimeWrapper_3_io_in = $signed(_T_517) < $signed(32'sh6); // @[package.scala 94:16:@33670.4]
  assign RetimeWrapper_4_clock = clock; // @[:@33677.4]
  assign RetimeWrapper_4_reset = reset; // @[:@33678.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33680.4]
  assign RetimeWrapper_4_io_in = $signed(_T_517) < $signed(32'sh3); // @[package.scala 94:16:@33679.4]
  assign RetimeWrapper_5_clock = clock; // @[:@33686.4]
  assign RetimeWrapper_5_reset = reset; // @[:@33687.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33689.4]
  assign RetimeWrapper_5_io_in = x429_sum_1_io_result; // @[package.scala 94:16:@33688.4]
  assign x436_sum_1_clock = clock; // @[:@33725.4]
  assign x436_sum_1_reset = reset; // @[:@33726.4]
  assign x436_sum_1_io_a = _T_574[31:0]; // @[Math.scala 151:17:@33727.4]
  assign x436_sum_1_io_b = _T_577[31:0]; // @[Math.scala 152:17:@33728.4]
  assign x436_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33729.4]
  assign x242_div_1_clock = clock; // @[:@33737.4]
  assign x242_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@33739.4]
  assign x242_div_1_io_flow = io_in_x202_TREADY; // @[Math.scala 330:20:@33741.4]
  assign RetimeWrapper_6_clock = clock; // @[:@33747.4]
  assign RetimeWrapper_6_reset = reset; // @[:@33748.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33750.4]
  assign RetimeWrapper_6_io_in = x436_sum_1_io_result; // @[package.scala 94:16:@33749.4]
  assign x243_sum_1_clock = clock; // @[:@33756.4]
  assign x243_sum_1_reset = reset; // @[:@33757.4]
  assign x243_sum_1_io_a = RetimeWrapper_6_io_out; // @[Math.scala 151:17:@33758.4]
  assign x243_sum_1_io_b = x242_div_1_io_result; // @[Math.scala 152:17:@33759.4]
  assign x243_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@33760.4]
  assign RetimeWrapper_7_clock = clock; // @[:@33766.4]
  assign RetimeWrapper_7_reset = reset; // @[:@33767.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33769.4]
  assign RetimeWrapper_7_io_in = $unsigned(_T_258); // @[package.scala 94:16:@33768.4]
  assign RetimeWrapper_8_clock = clock; // @[:@33775.4]
  assign RetimeWrapper_8_reset = reset; // @[:@33776.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33778.4]
  assign RetimeWrapper_8_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33777.4]
  assign RetimeWrapper_9_clock = clock; // @[:@33784.4]
  assign RetimeWrapper_9_reset = reset; // @[:@33785.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33787.4]
  assign RetimeWrapper_9_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@33786.4]
  assign RetimeWrapper_10_clock = clock; // @[:@33793.4]
  assign RetimeWrapper_10_reset = reset; // @[:@33794.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33796.4]
  assign RetimeWrapper_10_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33795.4]
  assign RetimeWrapper_11_clock = clock; // @[:@33802.4]
  assign RetimeWrapper_11_reset = reset; // @[:@33803.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33805.4]
  assign RetimeWrapper_11_io_in = x498_x430_D1 ? x499_x429_sum_D1_number : x432_sub_number; // @[package.scala 94:16:@33804.4]
  assign RetimeWrapper_12_clock = clock; // @[:@33813.4]
  assign RetimeWrapper_12_reset = reset; // @[:@33814.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33816.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33815.4]
  assign RetimeWrapper_13_clock = clock; // @[:@33834.4]
  assign RetimeWrapper_13_reset = reset; // @[:@33835.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33837.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@33836.4]
  assign RetimeWrapper_14_clock = clock; // @[:@33850.4]
  assign RetimeWrapper_14_reset = reset; // @[:@33851.4]
  assign RetimeWrapper_14_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@33853.4]
  assign RetimeWrapper_14_io_in = $signed(_T_633) < $signed(32'sh0); // @[package.scala 94:16:@33852.4]
  assign RetimeWrapper_15_clock = clock; // @[:@33859.4]
  assign RetimeWrapper_15_reset = reset; // @[:@33860.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33862.4]
  assign RetimeWrapper_15_io_in = __1_io_result; // @[package.scala 94:16:@33861.4]
  assign RetimeWrapper_16_clock = clock; // @[:@33873.4]
  assign RetimeWrapper_16_reset = reset; // @[:@33874.4]
  assign RetimeWrapper_16_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@33876.4]
  assign RetimeWrapper_16_io_in = $signed(_T_646) < $signed(32'sh0); // @[package.scala 94:16:@33875.4]
  assign RetimeWrapper_17_clock = clock; // @[:@33888.4]
  assign RetimeWrapper_17_reset = reset; // @[:@33889.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33891.4]
  assign RetimeWrapper_17_io_in = ~ x248; // @[package.scala 94:16:@33890.4]
  assign RetimeWrapper_18_clock = clock; // @[:@33897.4]
  assign RetimeWrapper_18_reset = reset; // @[:@33898.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33900.4]
  assign RetimeWrapper_18_io_in = $unsigned(_T_258); // @[package.scala 94:16:@33899.4]
  assign RetimeWrapper_19_clock = clock; // @[:@33906.4]
  assign RetimeWrapper_19_reset = reset; // @[:@33907.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33909.4]
  assign RetimeWrapper_19_io_in = x243_sum_1_io_result; // @[package.scala 94:16:@33908.4]
  assign RetimeWrapper_20_clock = clock; // @[:@33915.4]
  assign RetimeWrapper_20_reset = reset; // @[:@33916.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33918.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33917.4]
  assign RetimeWrapper_21_clock = clock; // @[:@33924.4]
  assign RetimeWrapper_21_reset = reset; // @[:@33925.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33927.4]
  assign RetimeWrapper_21_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33926.4]
  assign RetimeWrapper_22_clock = clock; // @[:@33933.4]
  assign RetimeWrapper_22_reset = reset; // @[:@33934.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33936.4]
  assign RetimeWrapper_22_io_in = x498_x430_D1 ? x499_x429_sum_D1_number : x432_sub_number; // @[package.scala 94:16:@33935.4]
  assign RetimeWrapper_23_clock = clock; // @[:@33945.4]
  assign RetimeWrapper_23_reset = reset; // @[:@33946.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33948.4]
  assign RetimeWrapper_23_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33947.4]
  assign x252_rdcol_1_clock = clock; // @[:@33968.4]
  assign x252_rdcol_1_reset = reset; // @[:@33969.4]
  assign x252_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@33970.4]
  assign x252_rdcol_1_io_b = 32'h1; // @[Math.scala 193:17:@33971.4]
  assign x252_rdcol_1_io_flow = io_in_x202_TREADY; // @[Math.scala 194:20:@33972.4]
  assign RetimeWrapper_24_clock = clock; // @[:@33983.4]
  assign RetimeWrapper_24_reset = reset; // @[:@33984.4]
  assign RetimeWrapper_24_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@33986.4]
  assign RetimeWrapper_24_io_in = $signed(_T_704) < $signed(32'sh0); // @[package.scala 94:16:@33985.4]
  assign RetimeWrapper_25_clock = clock; // @[:@33992.4]
  assign RetimeWrapper_25_reset = reset; // @[:@33993.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33995.4]
  assign RetimeWrapper_25_io_in = RetimeWrapper_14_io_out; // @[package.scala 94:16:@33994.4]
  assign x439_sum_1_clock = clock; // @[:@34035.4]
  assign x439_sum_1_reset = reset; // @[:@34036.4]
  assign x439_sum_1_io_a = _T_737 ? 32'h0 : _T_739; // @[Math.scala 151:17:@34037.4]
  assign x439_sum_1_io_b = $unsigned(_T_752); // @[Math.scala 152:17:@34038.4]
  assign x439_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34039.4]
  assign RetimeWrapper_26_clock = clock; // @[:@34058.4]
  assign RetimeWrapper_26_reset = reset; // @[:@34059.4]
  assign RetimeWrapper_26_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34061.4]
  assign RetimeWrapper_26_io_in = {_T_763,_T_764}; // @[package.scala 94:16:@34060.4]
  assign RetimeWrapper_27_clock = clock; // @[:@34076.4]
  assign RetimeWrapper_27_reset = reset; // @[:@34077.4]
  assign RetimeWrapper_27_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34080.4]
  assign RetimeWrapper_27_io_in = $unsigned(_T_795); // @[package.scala 94:16:@34079.4]
  assign x442_sum_1_clock = clock; // @[:@34089.4]
  assign x442_sum_1_reset = reset; // @[:@34090.4]
  assign x442_sum_1_io_a = _T_778 ? 32'h0 : _T_782; // @[Math.scala 151:17:@34091.4]
  assign x442_sum_1_io_b = $unsigned(_T_799); // @[Math.scala 152:17:@34092.4]
  assign x442_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34093.4]
  assign x445_sum_1_clock = clock; // @[:@34127.4]
  assign x445_sum_1_reset = reset; // @[:@34128.4]
  assign x445_sum_1_io_a = _T_825 ? 32'h0 : _T_827; // @[Math.scala 151:17:@34129.4]
  assign x445_sum_1_io_b = $unsigned(_T_840); // @[Math.scala 152:17:@34130.4]
  assign x445_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34131.4]
  assign x448_sum_1_clock = clock; // @[:@34165.4]
  assign x448_sum_1_reset = reset; // @[:@34166.4]
  assign x448_sum_1_io_a = _T_866 ? 32'h0 : _T_868; // @[Math.scala 151:17:@34167.4]
  assign x448_sum_1_io_b = $unsigned(_T_881); // @[Math.scala 152:17:@34168.4]
  assign x448_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34169.4]
  assign x451_sum_1_clock = clock; // @[:@34203.4]
  assign x451_sum_1_reset = reset; // @[:@34204.4]
  assign x451_sum_1_io_a = _T_907 ? 32'h0 : _T_909; // @[Math.scala 151:17:@34205.4]
  assign x451_sum_1_io_b = $unsigned(_T_922); // @[Math.scala 152:17:@34206.4]
  assign x451_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34207.4]
  assign x454_sum_1_clock = clock; // @[:@34241.4]
  assign x454_sum_1_reset = reset; // @[:@34242.4]
  assign x454_sum_1_io_a = _T_948 ? 32'h0 : _T_950; // @[Math.scala 151:17:@34243.4]
  assign x454_sum_1_io_b = $unsigned(_T_963); // @[Math.scala 152:17:@34244.4]
  assign x454_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34245.4]
  assign RetimeWrapper_28_clock = clock; // @[:@34256.4]
  assign RetimeWrapper_28_reset = reset; // @[:@34257.4]
  assign RetimeWrapper_28_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34259.4]
  assign RetimeWrapper_28_io_in = $signed(_T_973) < $signed(32'sh3); // @[package.scala 94:16:@34258.4]
  assign RetimeWrapper_29_clock = clock; // @[:@34270.4]
  assign RetimeWrapper_29_reset = reset; // @[:@34271.4]
  assign RetimeWrapper_29_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34273.4]
  assign RetimeWrapper_29_io_in = $signed(_T_973) < $signed(32'sh6); // @[package.scala 94:16:@34272.4]
  assign x457_sub_1_clock = clock; // @[:@34281.4]
  assign x457_sub_1_reset = reset; // @[:@34282.4]
  assign x457_sub_1_io_a = x454_sum_1_io_result; // @[Math.scala 192:17:@34283.4]
  assign x457_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@34284.4]
  assign x457_sub_1_io_flow = io_in_x202_TREADY; // @[Math.scala 194:20:@34285.4]
  assign RetimeWrapper_30_clock = clock; // @[:@34291.4]
  assign RetimeWrapper_30_reset = reset; // @[:@34292.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34294.4]
  assign RetimeWrapper_30_io_in = x454_sum_1_io_result; // @[package.scala 94:16:@34293.4]
  assign x257_div_1_clock = clock; // @[:@34305.4]
  assign x257_div_1_io_a = x252_rdcol_1_io_result; // @[Math.scala 328:17:@34307.4]
  assign x257_div_1_io_flow = io_in_x202_TREADY; // @[Math.scala 330:20:@34309.4]
  assign RetimeWrapper_31_clock = clock; // @[:@34315.4]
  assign RetimeWrapper_31_reset = reset; // @[:@34316.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34318.4]
  assign RetimeWrapper_31_io_in = x436_sum_1_io_result; // @[package.scala 94:16:@34317.4]
  assign x258_sum_1_clock = clock; // @[:@34324.4]
  assign x258_sum_1_reset = reset; // @[:@34325.4]
  assign x258_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@34326.4]
  assign x258_sum_1_io_b = x257_div_1_io_result; // @[Math.scala 152:17:@34327.4]
  assign x258_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34328.4]
  assign RetimeWrapper_32_clock = clock; // @[:@34334.4]
  assign RetimeWrapper_32_reset = reset; // @[:@34335.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34337.4]
  assign RetimeWrapper_32_io_in = ~ x254; // @[package.scala 94:16:@34336.4]
  assign RetimeWrapper_33_clock = clock; // @[:@34343.4]
  assign RetimeWrapper_33_reset = reset; // @[:@34344.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34346.4]
  assign RetimeWrapper_33_io_in = x455 ? x515_x454_sum_D1_number : x457_sub_number; // @[package.scala 94:16:@34345.4]
  assign RetimeWrapper_34_clock = clock; // @[:@34355.4]
  assign RetimeWrapper_34_reset = reset; // @[:@34356.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34358.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34357.4]
  assign x261_rdcol_1_clock = clock; // @[:@34378.4]
  assign x261_rdcol_1_reset = reset; // @[:@34379.4]
  assign x261_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@34380.4]
  assign x261_rdcol_1_io_b = 32'h2; // @[Math.scala 193:17:@34381.4]
  assign x261_rdcol_1_io_flow = io_in_x202_TREADY; // @[Math.scala 194:20:@34382.4]
  assign RetimeWrapper_35_clock = clock; // @[:@34395.4]
  assign RetimeWrapper_35_reset = reset; // @[:@34396.4]
  assign RetimeWrapper_35_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34398.4]
  assign RetimeWrapper_35_io_in = $signed(_T_1052) < $signed(32'sh0); // @[package.scala 94:16:@34397.4]
  assign x461_sum_1_clock = clock; // @[:@34438.4]
  assign x461_sum_1_reset = reset; // @[:@34439.4]
  assign x461_sum_1_io_a = _T_1082 ? 32'h0 : _T_1084; // @[Math.scala 151:17:@34440.4]
  assign x461_sum_1_io_b = $unsigned(_T_1097); // @[Math.scala 152:17:@34441.4]
  assign x461_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34442.4]
  assign RetimeWrapper_36_clock = clock; // @[:@34461.4]
  assign RetimeWrapper_36_reset = reset; // @[:@34462.4]
  assign RetimeWrapper_36_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34464.4]
  assign RetimeWrapper_36_io_in = {_T_1108,_T_1109}; // @[package.scala 94:16:@34463.4]
  assign RetimeWrapper_37_clock = clock; // @[:@34479.4]
  assign RetimeWrapper_37_reset = reset; // @[:@34480.4]
  assign RetimeWrapper_37_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34483.4]
  assign RetimeWrapper_37_io_in = $unsigned(_T_1140); // @[package.scala 94:16:@34482.4]
  assign x464_sum_1_clock = clock; // @[:@34492.4]
  assign x464_sum_1_reset = reset; // @[:@34493.4]
  assign x464_sum_1_io_a = _T_1123 ? 32'h0 : _T_1127; // @[Math.scala 151:17:@34494.4]
  assign x464_sum_1_io_b = $unsigned(_T_1144); // @[Math.scala 152:17:@34495.4]
  assign x464_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34496.4]
  assign x467_sum_1_clock = clock; // @[:@34530.4]
  assign x467_sum_1_reset = reset; // @[:@34531.4]
  assign x467_sum_1_io_a = _T_1170 ? 32'h0 : _T_1172; // @[Math.scala 151:17:@34532.4]
  assign x467_sum_1_io_b = $unsigned(_T_1185); // @[Math.scala 152:17:@34533.4]
  assign x467_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34534.4]
  assign x470_sum_1_clock = clock; // @[:@34568.4]
  assign x470_sum_1_reset = reset; // @[:@34569.4]
  assign x470_sum_1_io_a = _T_1211 ? 32'h0 : _T_1213; // @[Math.scala 151:17:@34570.4]
  assign x470_sum_1_io_b = $unsigned(_T_1226); // @[Math.scala 152:17:@34571.4]
  assign x470_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34572.4]
  assign x473_sum_1_clock = clock; // @[:@34606.4]
  assign x473_sum_1_reset = reset; // @[:@34607.4]
  assign x473_sum_1_io_a = _T_1252 ? 32'h0 : _T_1254; // @[Math.scala 151:17:@34608.4]
  assign x473_sum_1_io_b = $unsigned(_T_1267); // @[Math.scala 152:17:@34609.4]
  assign x473_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34610.4]
  assign x476_sum_1_clock = clock; // @[:@34644.4]
  assign x476_sum_1_reset = reset; // @[:@34645.4]
  assign x476_sum_1_io_a = _T_1293 ? 32'h0 : _T_1295; // @[Math.scala 151:17:@34646.4]
  assign x476_sum_1_io_b = $unsigned(_T_1308); // @[Math.scala 152:17:@34647.4]
  assign x476_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34648.4]
  assign RetimeWrapper_38_clock = clock; // @[:@34659.4]
  assign RetimeWrapper_38_reset = reset; // @[:@34660.4]
  assign RetimeWrapper_38_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34662.4]
  assign RetimeWrapper_38_io_in = $signed(_T_1318) < $signed(32'sh3); // @[package.scala 94:16:@34661.4]
  assign RetimeWrapper_39_clock = clock; // @[:@34673.4]
  assign RetimeWrapper_39_reset = reset; // @[:@34674.4]
  assign RetimeWrapper_39_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34676.4]
  assign RetimeWrapper_39_io_in = $signed(_T_1318) < $signed(32'sh6); // @[package.scala 94:16:@34675.4]
  assign x479_sub_1_clock = clock; // @[:@34684.4]
  assign x479_sub_1_reset = reset; // @[:@34685.4]
  assign x479_sub_1_io_a = x476_sum_1_io_result; // @[Math.scala 192:17:@34686.4]
  assign x479_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@34687.4]
  assign x479_sub_1_io_flow = io_in_x202_TREADY; // @[Math.scala 194:20:@34688.4]
  assign RetimeWrapper_40_clock = clock; // @[:@34694.4]
  assign RetimeWrapper_40_reset = reset; // @[:@34695.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34697.4]
  assign RetimeWrapper_40_io_in = x476_sum_1_io_result; // @[package.scala 94:16:@34696.4]
  assign x266_div_1_clock = clock; // @[:@34708.4]
  assign x266_div_1_io_a = x261_rdcol_1_io_result; // @[Math.scala 328:17:@34710.4]
  assign x266_div_1_io_flow = io_in_x202_TREADY; // @[Math.scala 330:20:@34712.4]
  assign x267_sum_1_clock = clock; // @[:@34718.4]
  assign x267_sum_1_reset = reset; // @[:@34719.4]
  assign x267_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@34720.4]
  assign x267_sum_1_io_b = x266_div_1_io_result; // @[Math.scala 152:17:@34721.4]
  assign x267_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34722.4]
  assign RetimeWrapper_41_clock = clock; // @[:@34728.4]
  assign RetimeWrapper_41_reset = reset; // @[:@34729.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34731.4]
  assign RetimeWrapper_41_io_in = x477 ? x519_x476_sum_D1_number : x479_sub_number; // @[package.scala 94:16:@34730.4]
  assign RetimeWrapper_42_clock = clock; // @[:@34737.4]
  assign RetimeWrapper_42_reset = reset; // @[:@34738.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34740.4]
  assign RetimeWrapper_42_io_in = ~ x263; // @[package.scala 94:16:@34739.4]
  assign RetimeWrapper_43_clock = clock; // @[:@34749.4]
  assign RetimeWrapper_43_reset = reset; // @[:@34750.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34752.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34751.4]
  assign x270_rdrow_1_clock = clock; // @[:@34772.4]
  assign x270_rdrow_1_reset = reset; // @[:@34773.4]
  assign x270_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@34774.4]
  assign x270_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@34775.4]
  assign x270_rdrow_1_io_flow = io_in_x202_TREADY; // @[Math.scala 194:20:@34776.4]
  assign RetimeWrapper_44_clock = clock; // @[:@34798.4]
  assign RetimeWrapper_44_reset = reset; // @[:@34799.4]
  assign RetimeWrapper_44_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34801.4]
  assign RetimeWrapper_44_io_in = $signed(_T_1394) < $signed(32'sh0); // @[package.scala 94:16:@34800.4]
  assign RetimeWrapper_45_clock = clock; // @[:@34807.4]
  assign RetimeWrapper_45_reset = reset; // @[:@34808.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34810.4]
  assign RetimeWrapper_45_io_in = RetimeWrapper_16_io_out; // @[package.scala 94:16:@34809.4]
  assign RetimeWrapper_46_clock = clock; // @[:@34829.4]
  assign RetimeWrapper_46_reset = reset; // @[:@34830.4]
  assign RetimeWrapper_46_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34833.4]
  assign RetimeWrapper_46_io_in = $unsigned(_T_1426); // @[package.scala 94:16:@34832.4]
  assign RetimeWrapper_47_clock = clock; // @[:@34855.4]
  assign RetimeWrapper_47_reset = reset; // @[:@34856.4]
  assign RetimeWrapper_47_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@34858.4]
  assign RetimeWrapper_47_io_in = {_T_1438,_T_1439}; // @[package.scala 94:16:@34857.4]
  assign x485_sum_1_clock = clock; // @[:@34876.4]
  assign x485_sum_1_reset = reset; // @[:@34877.4]
  assign x485_sum_1_io_a = _T_1462[31:0]; // @[Math.scala 151:17:@34878.4]
  assign x485_sum_1_io_b = _T_1465[31:0]; // @[Math.scala 152:17:@34879.4]
  assign x485_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34880.4]
  assign RetimeWrapper_48_clock = clock; // @[:@34886.4]
  assign RetimeWrapper_48_reset = reset; // @[:@34887.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34889.4]
  assign RetimeWrapper_48_io_in = x242_div_1_io_result; // @[package.scala 94:16:@34888.4]
  assign RetimeWrapper_49_clock = clock; // @[:@34895.4]
  assign RetimeWrapper_49_reset = reset; // @[:@34896.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34898.4]
  assign RetimeWrapper_49_io_in = x485_sum_1_io_result; // @[package.scala 94:16:@34897.4]
  assign x278_sum_1_clock = clock; // @[:@34904.4]
  assign x278_sum_1_reset = reset; // @[:@34905.4]
  assign x278_sum_1_io_a = RetimeWrapper_49_io_out; // @[Math.scala 151:17:@34906.4]
  assign x278_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@34907.4]
  assign x278_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34908.4]
  assign RetimeWrapper_50_clock = clock; // @[:@34914.4]
  assign RetimeWrapper_50_reset = reset; // @[:@34915.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34917.4]
  assign RetimeWrapper_50_io_in = ~ x273; // @[package.scala 94:16:@34916.4]
  assign RetimeWrapper_51_clock = clock; // @[:@34923.4]
  assign RetimeWrapper_51_reset = reset; // @[:@34924.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34926.4]
  assign RetimeWrapper_51_io_in = x278_sum_1_io_result; // @[package.scala 94:16:@34925.4]
  assign RetimeWrapper_52_clock = clock; // @[:@34932.4]
  assign RetimeWrapper_52_reset = reset; // @[:@34933.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34935.4]
  assign RetimeWrapper_52_io_in = $unsigned(_T_1430); // @[package.scala 94:16:@34934.4]
  assign RetimeWrapper_53_clock = clock; // @[:@34944.4]
  assign RetimeWrapper_53_reset = reset; // @[:@34945.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34947.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34946.4]
  assign RetimeWrapper_54_clock = clock; // @[:@34971.4]
  assign RetimeWrapper_54_reset = reset; // @[:@34972.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34974.4]
  assign RetimeWrapper_54_io_in = x485_sum_1_io_result; // @[package.scala 94:16:@34973.4]
  assign x283_sum_1_clock = clock; // @[:@34982.4]
  assign x283_sum_1_reset = reset; // @[:@34983.4]
  assign x283_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@34984.4]
  assign x283_sum_1_io_b = x257_div_1_io_result; // @[Math.scala 152:17:@34985.4]
  assign x283_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@34986.4]
  assign RetimeWrapper_55_clock = clock; // @[:@34992.4]
  assign RetimeWrapper_55_reset = reset; // @[:@34993.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34995.4]
  assign RetimeWrapper_55_io_in = ~ x281; // @[package.scala 94:16:@34994.4]
  assign RetimeWrapper_56_clock = clock; // @[:@35004.4]
  assign RetimeWrapper_56_reset = reset; // @[:@35005.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35007.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35006.4]
  assign x288_sum_1_clock = clock; // @[:@35031.4]
  assign x288_sum_1_reset = reset; // @[:@35032.4]
  assign x288_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@35033.4]
  assign x288_sum_1_io_b = x266_div_1_io_result; // @[Math.scala 152:17:@35034.4]
  assign x288_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35035.4]
  assign RetimeWrapper_57_clock = clock; // @[:@35041.4]
  assign RetimeWrapper_57_reset = reset; // @[:@35042.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35044.4]
  assign RetimeWrapper_57_io_in = ~ x286; // @[package.scala 94:16:@35043.4]
  assign RetimeWrapper_58_clock = clock; // @[:@35053.4]
  assign RetimeWrapper_58_reset = reset; // @[:@35054.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35056.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35055.4]
  assign x291_rdrow_1_clock = clock; // @[:@35076.4]
  assign x291_rdrow_1_reset = reset; // @[:@35077.4]
  assign x291_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@35078.4]
  assign x291_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@35079.4]
  assign x291_rdrow_1_io_flow = io_in_x202_TREADY; // @[Math.scala 194:20:@35080.4]
  assign RetimeWrapper_59_clock = clock; // @[:@35102.4]
  assign RetimeWrapper_59_reset = reset; // @[:@35103.4]
  assign RetimeWrapper_59_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@35105.4]
  assign RetimeWrapper_59_io_in = $signed(_T_1583) < $signed(32'sh0); // @[package.scala 94:16:@35104.4]
  assign RetimeWrapper_60_clock = clock; // @[:@35124.4]
  assign RetimeWrapper_60_reset = reset; // @[:@35125.4]
  assign RetimeWrapper_60_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@35128.4]
  assign RetimeWrapper_60_io_in = $unsigned(_T_1612); // @[package.scala 94:16:@35127.4]
  assign RetimeWrapper_61_clock = clock; // @[:@35150.4]
  assign RetimeWrapper_61_reset = reset; // @[:@35151.4]
  assign RetimeWrapper_61_io_flow = io_in_x202_TREADY; // @[package.scala 95:18:@35153.4]
  assign RetimeWrapper_61_io_in = {_T_1624,_T_1625}; // @[package.scala 94:16:@35152.4]
  assign x490_sum_1_clock = clock; // @[:@35171.4]
  assign x490_sum_1_reset = reset; // @[:@35172.4]
  assign x490_sum_1_io_a = _T_1648[31:0]; // @[Math.scala 151:17:@35173.4]
  assign x490_sum_1_io_b = _T_1651[31:0]; // @[Math.scala 152:17:@35174.4]
  assign x490_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35175.4]
  assign RetimeWrapper_62_clock = clock; // @[:@35181.4]
  assign RetimeWrapper_62_reset = reset; // @[:@35182.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35184.4]
  assign RetimeWrapper_62_io_in = x490_sum_1_io_result; // @[package.scala 94:16:@35183.4]
  assign x299_sum_1_clock = clock; // @[:@35190.4]
  assign x299_sum_1_reset = reset; // @[:@35191.4]
  assign x299_sum_1_io_a = RetimeWrapper_62_io_out; // @[Math.scala 151:17:@35192.4]
  assign x299_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@35193.4]
  assign x299_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35194.4]
  assign RetimeWrapper_63_clock = clock; // @[:@35200.4]
  assign RetimeWrapper_63_reset = reset; // @[:@35201.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35203.4]
  assign RetimeWrapper_63_io_in = x299_sum_1_io_result; // @[package.scala 94:16:@35202.4]
  assign RetimeWrapper_64_clock = clock; // @[:@35209.4]
  assign RetimeWrapper_64_reset = reset; // @[:@35210.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35212.4]
  assign RetimeWrapper_64_io_in = $unsigned(_T_1616); // @[package.scala 94:16:@35211.4]
  assign RetimeWrapper_65_clock = clock; // @[:@35218.4]
  assign RetimeWrapper_65_reset = reset; // @[:@35219.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35221.4]
  assign RetimeWrapper_65_io_in = ~ x294; // @[package.scala 94:16:@35220.4]
  assign RetimeWrapper_66_clock = clock; // @[:@35230.4]
  assign RetimeWrapper_66_reset = reset; // @[:@35231.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35233.4]
  assign RetimeWrapper_66_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35232.4]
  assign RetimeWrapper_67_clock = clock; // @[:@35257.4]
  assign RetimeWrapper_67_reset = reset; // @[:@35258.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35260.4]
  assign RetimeWrapper_67_io_in = x490_sum_1_io_result; // @[package.scala 94:16:@35259.4]
  assign x304_sum_1_clock = clock; // @[:@35266.4]
  assign x304_sum_1_reset = reset; // @[:@35267.4]
  assign x304_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@35268.4]
  assign x304_sum_1_io_b = x257_div_1_io_result; // @[Math.scala 152:17:@35269.4]
  assign x304_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35270.4]
  assign RetimeWrapper_68_clock = clock; // @[:@35276.4]
  assign RetimeWrapper_68_reset = reset; // @[:@35277.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35279.4]
  assign RetimeWrapper_68_io_in = ~ x302; // @[package.scala 94:16:@35278.4]
  assign RetimeWrapper_69_clock = clock; // @[:@35288.4]
  assign RetimeWrapper_69_reset = reset; // @[:@35289.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35291.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35290.4]
  assign x309_sum_1_clock = clock; // @[:@35315.4]
  assign x309_sum_1_reset = reset; // @[:@35316.4]
  assign x309_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@35317.4]
  assign x309_sum_1_io_b = x266_div_1_io_result; // @[Math.scala 152:17:@35318.4]
  assign x309_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35319.4]
  assign RetimeWrapper_70_clock = clock; // @[:@35325.4]
  assign RetimeWrapper_70_reset = reset; // @[:@35326.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35328.4]
  assign RetimeWrapper_70_io_in = ~ x307; // @[package.scala 94:16:@35327.4]
  assign RetimeWrapper_71_clock = clock; // @[:@35337.4]
  assign RetimeWrapper_71_reset = reset; // @[:@35338.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35340.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35339.4]
  assign x312_1_clock = clock; // @[:@35360.4]
  assign x312_1_io_a = x233_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@35362.4]
  assign x312_1_io_b = 32'h1; // @[Math.scala 264:17:@35363.4]
  assign x312_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35364.4]
  assign x313_1_clock = clock; // @[:@35372.4]
  assign x313_1_io_a = x233_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@35374.4]
  assign x313_1_io_b = 32'h2; // @[Math.scala 264:17:@35375.4]
  assign x313_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35376.4]
  assign x314_1_clock = clock; // @[:@35384.4]
  assign x314_1_io_a = x233_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@35386.4]
  assign x314_1_io_b = 32'h1; // @[Math.scala 264:17:@35387.4]
  assign x314_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35388.4]
  assign x315_1_clock = clock; // @[:@35396.4]
  assign x315_1_io_a = x233_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@35398.4]
  assign x315_1_io_b = 32'h2; // @[Math.scala 264:17:@35399.4]
  assign x315_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35400.4]
  assign x316_1_clock = clock; // @[:@35410.4]
  assign x316_1_io_a = x233_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@35412.4]
  assign x316_1_io_b = 32'h4; // @[Math.scala 264:17:@35413.4]
  assign x316_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35414.4]
  assign x317_1_clock = clock; // @[:@35422.4]
  assign x317_1_io_a = x233_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@35424.4]
  assign x317_1_io_b = 32'h2; // @[Math.scala 264:17:@35425.4]
  assign x317_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35426.4]
  assign x318_1_clock = clock; // @[:@35434.4]
  assign x318_1_io_a = x233_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@35436.4]
  assign x318_1_io_b = 32'h1; // @[Math.scala 264:17:@35437.4]
  assign x318_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35438.4]
  assign x319_1_clock = clock; // @[:@35446.4]
  assign x319_1_io_a = x233_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@35448.4]
  assign x319_1_io_b = 32'h2; // @[Math.scala 264:17:@35449.4]
  assign x319_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35450.4]
  assign x320_1_clock = clock; // @[:@35458.4]
  assign x320_1_io_a = x233_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@35460.4]
  assign x320_1_io_b = 32'h1; // @[Math.scala 264:17:@35461.4]
  assign x320_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35462.4]
  assign x321_x7_1_clock = clock; // @[:@35468.4]
  assign x321_x7_1_reset = reset; // @[:@35469.4]
  assign x321_x7_1_io_a = x312_1_io_result; // @[Math.scala 151:17:@35470.4]
  assign x321_x7_1_io_b = x313_1_io_result; // @[Math.scala 152:17:@35471.4]
  assign x321_x7_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35472.4]
  assign x322_x8_1_clock = clock; // @[:@35478.4]
  assign x322_x8_1_reset = reset; // @[:@35479.4]
  assign x322_x8_1_io_a = x314_1_io_result; // @[Math.scala 151:17:@35480.4]
  assign x322_x8_1_io_b = x315_1_io_result; // @[Math.scala 152:17:@35481.4]
  assign x322_x8_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35482.4]
  assign x323_x7_1_clock = clock; // @[:@35488.4]
  assign x323_x7_1_reset = reset; // @[:@35489.4]
  assign x323_x7_1_io_a = x316_1_io_result; // @[Math.scala 151:17:@35490.4]
  assign x323_x7_1_io_b = x317_1_io_result; // @[Math.scala 152:17:@35491.4]
  assign x323_x7_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35492.4]
  assign x324_x8_1_clock = clock; // @[:@35498.4]
  assign x324_x8_1_reset = reset; // @[:@35499.4]
  assign x324_x8_1_io_a = x318_1_io_result; // @[Math.scala 151:17:@35500.4]
  assign x324_x8_1_io_b = x319_1_io_result; // @[Math.scala 152:17:@35501.4]
  assign x324_x8_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35502.4]
  assign x325_x7_1_clock = clock; // @[:@35508.4]
  assign x325_x7_1_reset = reset; // @[:@35509.4]
  assign x325_x7_1_io_a = x321_x7_1_io_result; // @[Math.scala 151:17:@35510.4]
  assign x325_x7_1_io_b = x322_x8_1_io_result; // @[Math.scala 152:17:@35511.4]
  assign x325_x7_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35512.4]
  assign x326_x8_1_clock = clock; // @[:@35518.4]
  assign x326_x8_1_reset = reset; // @[:@35519.4]
  assign x326_x8_1_io_a = x323_x7_1_io_result; // @[Math.scala 151:17:@35520.4]
  assign x326_x8_1_io_b = x324_x8_1_io_result; // @[Math.scala 152:17:@35521.4]
  assign x326_x8_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35522.4]
  assign x327_x7_1_clock = clock; // @[:@35528.4]
  assign x327_x7_1_reset = reset; // @[:@35529.4]
  assign x327_x7_1_io_a = x325_x7_1_io_result; // @[Math.scala 151:17:@35530.4]
  assign x327_x7_1_io_b = x326_x8_1_io_result; // @[Math.scala 152:17:@35531.4]
  assign x327_x7_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35532.4]
  assign RetimeWrapper_72_clock = clock; // @[:@35538.4]
  assign RetimeWrapper_72_reset = reset; // @[:@35539.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35541.4]
  assign RetimeWrapper_72_io_in = x320_1_io_result; // @[package.scala 94:16:@35540.4]
  assign x328_sum_1_clock = clock; // @[:@35547.4]
  assign x328_sum_1_reset = reset; // @[:@35548.4]
  assign x328_sum_1_io_a = x327_x7_1_io_result; // @[Math.scala 151:17:@35549.4]
  assign x328_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@35550.4]
  assign x328_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35551.4]
  assign x329_1_io_b = x328_sum_1_io_result; // @[Math.scala 721:17:@35559.4]
  assign x330_mul_1_clock = clock; // @[:@35568.4]
  assign x330_mul_1_io_a = x329_1_io_result; // @[Math.scala 263:17:@35570.4]
  assign x330_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@35571.4]
  assign x330_mul_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35572.4]
  assign x331_1_io_b = x330_mul_1_io_result; // @[Math.scala 721:17:@35580.4]
  assign RetimeWrapper_73_clock = clock; // @[:@35587.4]
  assign RetimeWrapper_73_reset = reset; // @[:@35588.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35590.4]
  assign RetimeWrapper_73_io_in = $unsigned(_T_258); // @[package.scala 94:16:@35589.4]
  assign RetimeWrapper_74_clock = clock; // @[:@35596.4]
  assign RetimeWrapper_74_reset = reset; // @[:@35597.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35599.4]
  assign RetimeWrapper_74_io_in = x243_sum_1_io_result; // @[package.scala 94:16:@35598.4]
  assign RetimeWrapper_75_clock = clock; // @[:@35605.4]
  assign RetimeWrapper_75_reset = reset; // @[:@35606.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35608.4]
  assign RetimeWrapper_75_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@35607.4]
  assign RetimeWrapper_76_clock = clock; // @[:@35614.4]
  assign RetimeWrapper_76_reset = reset; // @[:@35615.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35617.4]
  assign RetimeWrapper_76_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@35616.4]
  assign RetimeWrapper_77_clock = clock; // @[:@35623.4]
  assign RetimeWrapper_77_reset = reset; // @[:@35624.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35626.4]
  assign RetimeWrapper_77_io_in = x331_1_io_result; // @[package.scala 94:16:@35625.4]
  assign RetimeWrapper_78_clock = clock; // @[:@35632.4]
  assign RetimeWrapper_78_reset = reset; // @[:@35633.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35635.4]
  assign RetimeWrapper_78_io_in = x498_x430_D1 ? x499_x429_sum_D1_number : x432_sub_number; // @[package.scala 94:16:@35634.4]
  assign RetimeWrapper_79_clock = clock; // @[:@35643.4]
  assign RetimeWrapper_79_reset = reset; // @[:@35644.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35646.4]
  assign RetimeWrapper_79_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35645.4]
  assign RetimeWrapper_80_clock = clock; // @[:@35664.4]
  assign RetimeWrapper_80_reset = reset; // @[:@35665.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35667.4]
  assign RetimeWrapper_80_io_in = ~ x248; // @[package.scala 94:16:@35666.4]
  assign RetimeWrapper_81_clock = clock; // @[:@35673.4]
  assign RetimeWrapper_81_reset = reset; // @[:@35674.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35676.4]
  assign RetimeWrapper_81_io_in = $unsigned(_T_258); // @[package.scala 94:16:@35675.4]
  assign RetimeWrapper_82_clock = clock; // @[:@35682.4]
  assign RetimeWrapper_82_reset = reset; // @[:@35683.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35685.4]
  assign RetimeWrapper_82_io_in = x243_sum_1_io_result; // @[package.scala 94:16:@35684.4]
  assign RetimeWrapper_83_clock = clock; // @[:@35691.4]
  assign RetimeWrapper_83_reset = reset; // @[:@35692.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35694.4]
  assign RetimeWrapper_83_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@35693.4]
  assign RetimeWrapper_84_clock = clock; // @[:@35700.4]
  assign RetimeWrapper_84_reset = reset; // @[:@35701.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35703.4]
  assign RetimeWrapper_84_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@35702.4]
  assign RetimeWrapper_85_clock = clock; // @[:@35709.4]
  assign RetimeWrapper_85_reset = reset; // @[:@35710.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35712.4]
  assign RetimeWrapper_85_io_in = x498_x430_D1 ? x499_x429_sum_D1_number : x432_sub_number; // @[package.scala 94:16:@35711.4]
  assign RetimeWrapper_86_clock = clock; // @[:@35721.4]
  assign RetimeWrapper_86_reset = reset; // @[:@35722.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35724.4]
  assign RetimeWrapper_86_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35723.4]
  assign RetimeWrapper_87_clock = clock; // @[:@35742.4]
  assign RetimeWrapper_87_reset = reset; // @[:@35743.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35745.4]
  assign RetimeWrapper_87_io_in = ~ x254; // @[package.scala 94:16:@35744.4]
  assign RetimeWrapper_88_clock = clock; // @[:@35751.4]
  assign RetimeWrapper_88_reset = reset; // @[:@35752.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35754.4]
  assign RetimeWrapper_88_io_in = x455 ? x515_x454_sum_D1_number : x457_sub_number; // @[package.scala 94:16:@35753.4]
  assign RetimeWrapper_89_clock = clock; // @[:@35760.4]
  assign RetimeWrapper_89_reset = reset; // @[:@35761.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35763.4]
  assign RetimeWrapper_89_io_in = x258_sum_1_io_result; // @[package.scala 94:16:@35762.4]
  assign RetimeWrapper_90_clock = clock; // @[:@35772.4]
  assign RetimeWrapper_90_reset = reset; // @[:@35773.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35775.4]
  assign RetimeWrapper_90_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35774.4]
  assign RetimeWrapper_91_clock = clock; // @[:@35793.4]
  assign RetimeWrapper_91_reset = reset; // @[:@35794.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35796.4]
  assign RetimeWrapper_91_io_in = ~ x273; // @[package.scala 94:16:@35795.4]
  assign RetimeWrapper_92_clock = clock; // @[:@35802.4]
  assign RetimeWrapper_92_reset = reset; // @[:@35803.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35805.4]
  assign RetimeWrapper_92_io_in = x278_sum_1_io_result; // @[package.scala 94:16:@35804.4]
  assign RetimeWrapper_93_clock = clock; // @[:@35811.4]
  assign RetimeWrapper_93_reset = reset; // @[:@35812.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35814.4]
  assign RetimeWrapper_93_io_in = $unsigned(_T_1430); // @[package.scala 94:16:@35813.4]
  assign RetimeWrapper_94_clock = clock; // @[:@35823.4]
  assign RetimeWrapper_94_reset = reset; // @[:@35824.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35826.4]
  assign RetimeWrapper_94_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35825.4]
  assign RetimeWrapper_95_clock = clock; // @[:@35844.4]
  assign RetimeWrapper_95_reset = reset; // @[:@35845.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35847.4]
  assign RetimeWrapper_95_io_in = ~ x281; // @[package.scala 94:16:@35846.4]
  assign RetimeWrapper_96_clock = clock; // @[:@35853.4]
  assign RetimeWrapper_96_reset = reset; // @[:@35854.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35856.4]
  assign RetimeWrapper_96_io_in = x283_sum_1_io_result; // @[package.scala 94:16:@35855.4]
  assign RetimeWrapper_97_clock = clock; // @[:@35865.4]
  assign RetimeWrapper_97_reset = reset; // @[:@35866.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35868.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35867.4]
  assign x343_1_clock = clock; // @[:@35888.4]
  assign x343_1_io_a = x234_lb2_0_io_rPort_0_output_0; // @[Math.scala 263:17:@35890.4]
  assign x343_1_io_b = 32'h1; // @[Math.scala 264:17:@35891.4]
  assign x343_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35892.4]
  assign x344_1_clock = clock; // @[:@35902.4]
  assign x344_1_io_a = x234_lb2_0_io_rPort_1_output_0; // @[Math.scala 263:17:@35904.4]
  assign x344_1_io_b = 32'h2; // @[Math.scala 264:17:@35905.4]
  assign x344_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35906.4]
  assign x345_1_clock = clock; // @[:@35914.4]
  assign x345_1_io_a = x234_lb2_0_io_rPort_2_output_0; // @[Math.scala 263:17:@35916.4]
  assign x345_1_io_b = 32'h4; // @[Math.scala 264:17:@35917.4]
  assign x345_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35918.4]
  assign x346_1_clock = clock; // @[:@35926.4]
  assign x346_1_io_a = x234_lb2_0_io_rPort_3_output_0; // @[Math.scala 263:17:@35928.4]
  assign x346_1_io_b = 32'h1; // @[Math.scala 264:17:@35929.4]
  assign x346_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35930.4]
  assign x347_x9_1_clock = clock; // @[:@35936.4]
  assign x347_x9_1_reset = reset; // @[:@35937.4]
  assign x347_x9_1_io_a = x343_1_io_result; // @[Math.scala 151:17:@35938.4]
  assign x347_x9_1_io_b = x344_1_io_result; // @[Math.scala 152:17:@35939.4]
  assign x347_x9_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35940.4]
  assign x348_x10_1_clock = clock; // @[:@35946.4]
  assign x348_x10_1_reset = reset; // @[:@35947.4]
  assign x348_x10_1_io_a = x345_1_io_result; // @[Math.scala 151:17:@35948.4]
  assign x348_x10_1_io_b = x346_1_io_result; // @[Math.scala 152:17:@35949.4]
  assign x348_x10_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35950.4]
  assign x349_sum_1_clock = clock; // @[:@35956.4]
  assign x349_sum_1_reset = reset; // @[:@35957.4]
  assign x349_sum_1_io_a = x347_x9_1_io_result; // @[Math.scala 151:17:@35958.4]
  assign x349_sum_1_io_b = x348_x10_1_io_result; // @[Math.scala 152:17:@35959.4]
  assign x349_sum_1_io_flow = io_in_x202_TREADY; // @[Math.scala 153:20:@35960.4]
  assign x350_1_io_b = x349_sum_1_io_result; // @[Math.scala 721:17:@35968.4]
  assign x351_mul_1_clock = clock; // @[:@35977.4]
  assign x351_mul_1_io_a = x350_1_io_result; // @[Math.scala 263:17:@35979.4]
  assign x351_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@35980.4]
  assign x351_mul_1_io_flow = io_in_x202_TREADY; // @[Math.scala 265:20:@35981.4]
  assign x352_1_io_b = x351_mul_1_io_result; // @[Math.scala 721:17:@35989.4]
  assign RetimeWrapper_98_clock = clock; // @[:@36000.4]
  assign RetimeWrapper_98_reset = reset; // @[:@36001.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36003.4]
  assign RetimeWrapper_98_io_in = x352_1_io_result; // @[package.scala 94:16:@36002.4]
  assign RetimeWrapper_99_clock = clock; // @[:@36009.4]
  assign RetimeWrapper_99_reset = reset; // @[:@36010.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36012.4]
  assign RetimeWrapper_99_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@36011.4]
  assign RetimeWrapper_100_clock = clock; // @[:@36018.4]
  assign RetimeWrapper_100_reset = reset; // @[:@36019.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36021.4]
  assign RetimeWrapper_100_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@36020.4]
  assign RetimeWrapper_101_clock = clock; // @[:@36027.4]
  assign RetimeWrapper_101_reset = reset; // @[:@36028.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36030.4]
  assign RetimeWrapper_101_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@36029.4]
endmodule
module x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1( // @[:@36048.2]
  input          clock, // @[:@36049.4]
  input          reset, // @[:@36050.4]
  output         io_in_x202_TVALID, // @[:@36051.4]
  input          io_in_x202_TREADY, // @[:@36051.4]
  output [255:0] io_in_x202_TDATA, // @[:@36051.4]
  input          io_in_x201_TVALID, // @[:@36051.4]
  output         io_in_x201_TREADY, // @[:@36051.4]
  input  [255:0] io_in_x201_TDATA, // @[:@36051.4]
  input  [7:0]   io_in_x201_TID, // @[:@36051.4]
  input  [7:0]   io_in_x201_TDEST, // @[:@36051.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@36051.4]
  input          io_sigsIn_smChildAcks_0, // @[:@36051.4]
  output         io_sigsOut_smDoneIn_0, // @[:@36051.4]
  input          io_rr // @[:@36051.4]
);
  wire  x226_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire  x226_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire  x226_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire  x226_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire [12:0] x226_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire [12:0] x226_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire  x226_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire  x226_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire  x226_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@36085.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36173.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36173.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36173.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36173.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36173.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36215.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36215.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36215.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36215.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36215.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@36223.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@36223.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@36223.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@36223.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@36223.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TVALID; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TREADY; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire [255:0] x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TDATA; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TREADY; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire [255:0] x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TDATA; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire [7:0] x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TID; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire [7:0] x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TDEST; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire [31:0] x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire [31:0] x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
  wire  _T_240; // @[package.scala 96:25:@36178.4 package.scala 96:25:@36179.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x358_outr_UnitPipe.scala 69:66:@36184.4]
  wire  _T_253; // @[package.scala 96:25:@36220.4 package.scala 96:25:@36221.4]
  wire  _T_259; // @[package.scala 96:25:@36228.4 package.scala 96:25:@36229.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@36231.4]
  wire  x357_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@36232.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@36240.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@36241.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@36253.4]
  x209_ctrchain x226_ctrchain ( // @[SpatialBlocks.scala 37:22:@36085.4]
    .clock(x226_ctrchain_clock),
    .reset(x226_ctrchain_reset),
    .io_input_reset(x226_ctrchain_io_input_reset),
    .io_input_enable(x226_ctrchain_io_input_enable),
    .io_output_counts_1(x226_ctrchain_io_output_counts_1),
    .io_output_counts_0(x226_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x226_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x226_ctrchain_io_output_oobs_1),
    .io_output_done(x226_ctrchain_io_output_done)
  );
  x357_inr_Foreach_SAMPLER_BOX_sm x357_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 32:18:@36145.4]
    .clock(x357_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x357_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x357_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x357_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x357_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x357_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x357_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x357_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x357_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36173.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36215.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@36223.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1 x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 680:24:@36257.4]
    .clock(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x202_TVALID(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TVALID),
    .io_in_x202_TREADY(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TREADY),
    .io_in_x202_TDATA(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TDATA),
    .io_in_x201_TREADY(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TREADY),
    .io_in_x201_TDATA(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TDATA),
    .io_in_x201_TID(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TID),
    .io_in_x201_TDEST(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TDEST),
    .io_sigsIn_backpressure(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@36178.4 package.scala 96:25:@36179.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x201_TVALID | x357_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x358_outr_UnitPipe.scala 69:66:@36184.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36220.4 package.scala 96:25:@36221.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@36228.4 package.scala 96:25:@36229.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@36231.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@36232.4]
  assign _T_264 = x357_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@36240.4]
  assign _T_265 = ~ x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@36241.4]
  assign _T_272 = x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@36253.4]
  assign io_in_x202_TVALID = x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TVALID; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 48:23:@36316.4]
  assign io_in_x202_TDATA = x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TDATA; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 48:23:@36314.4]
  assign io_in_x201_TREADY = x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TREADY; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 49:23:@36324.4]
  assign io_sigsOut_smDoneIn_0 = x357_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@36238.4]
  assign x226_ctrchain_clock = clock; // @[:@36086.4]
  assign x226_ctrchain_reset = reset; // @[:@36087.4]
  assign x226_ctrchain_io_input_reset = x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@36256.4]
  assign x226_ctrchain_io_input_enable = _T_272 & x357_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@36208.4 SpatialBlocks.scala 159:42:@36255.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@36146.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@36147.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sm_io_enable = x357_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x357_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@36235.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x358_outr_UnitPipe.scala 67:50:@36181.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@36237.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x202_TREADY | x357_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@36209.4]
  assign x357_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x358_outr_UnitPipe.scala 71:48:@36187.4]
  assign RetimeWrapper_clock = clock; // @[:@36174.4]
  assign RetimeWrapper_reset = reset; // @[:@36175.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36177.4]
  assign RetimeWrapper_io_in = x226_ctrchain_io_output_done; // @[package.scala 94:16:@36176.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36216.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36217.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36219.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@36218.4]
  assign RetimeWrapper_2_clock = clock; // @[:@36224.4]
  assign RetimeWrapper_2_reset = reset; // @[:@36225.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@36227.4]
  assign RetimeWrapper_2_io_in = x357_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@36226.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@36258.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@36259.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x202_TREADY = io_in_x202_TREADY; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 48:23:@36315.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TDATA = io_in_x201_TDATA; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 49:23:@36323.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TID = io_in_x201_TID; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 49:23:@36319.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x201_TDEST = io_in_x201_TDEST; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 49:23:@36318.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x202_TREADY | x357_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 685:22:@36342.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 685:22:@36340.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x357_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 685:22:@36338.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x226_ctrchain_io_output_counts_1[12]}},x226_ctrchain_io_output_counts_1}; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 685:22:@36333.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x226_ctrchain_io_output_counts_0[12]}},x226_ctrchain_io_output_counts_0}; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 685:22:@36332.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x226_ctrchain_io_output_oobs_0; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 685:22:@36330.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x226_ctrchain_io_output_oobs_1; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 685:22:@36331.4]
  assign x357_inr_Foreach_SAMPLER_BOX_kernelx357_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x357_inr_Foreach_SAMPLER_BOX.scala 684:18:@36326.4]
endmodule
module x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1( // @[:@36356.2]
  input          clock, // @[:@36357.4]
  input          reset, // @[:@36358.4]
  output         io_in_x202_TVALID, // @[:@36359.4]
  input          io_in_x202_TREADY, // @[:@36359.4]
  output [255:0] io_in_x202_TDATA, // @[:@36359.4]
  input          io_in_x201_TVALID, // @[:@36359.4]
  output         io_in_x201_TREADY, // @[:@36359.4]
  input  [255:0] io_in_x201_TDATA, // @[:@36359.4]
  input  [7:0]   io_in_x201_TID, // @[:@36359.4]
  input  [7:0]   io_in_x201_TDEST, // @[:@36359.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@36359.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@36359.4]
  input          io_sigsIn_smChildAcks_0, // @[:@36359.4]
  input          io_sigsIn_smChildAcks_1, // @[:@36359.4]
  output         io_sigsOut_smDoneIn_0, // @[:@36359.4]
  output         io_sigsOut_smDoneIn_1, // @[:@36359.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@36359.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@36359.4]
  input          io_rr // @[:@36359.4]
);
  wire  x204_fifoinraw_0_clock; // @[m_x204_fifoinraw_0.scala 27:17:@36373.4]
  wire  x204_fifoinraw_0_reset; // @[m_x204_fifoinraw_0.scala 27:17:@36373.4]
  wire  x205_fifoinpacked_0_clock; // @[m_x205_fifoinpacked_0.scala 27:17:@36397.4]
  wire  x205_fifoinpacked_0_reset; // @[m_x205_fifoinpacked_0.scala 27:17:@36397.4]
  wire  x205_fifoinpacked_0_io_wPort_0_en_0; // @[m_x205_fifoinpacked_0.scala 27:17:@36397.4]
  wire  x205_fifoinpacked_0_io_full; // @[m_x205_fifoinpacked_0.scala 27:17:@36397.4]
  wire  x205_fifoinpacked_0_io_active_0_in; // @[m_x205_fifoinpacked_0.scala 27:17:@36397.4]
  wire  x205_fifoinpacked_0_io_active_0_out; // @[m_x205_fifoinpacked_0.scala 27:17:@36397.4]
  wire  x206_fifooutraw_0_clock; // @[m_x206_fifooutraw_0.scala 27:17:@36421.4]
  wire  x206_fifooutraw_0_reset; // @[m_x206_fifooutraw_0.scala 27:17:@36421.4]
  wire  x209_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire  x209_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire  x209_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire  x209_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire [12:0] x209_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire [12:0] x209_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire  x209_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire  x209_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire  x209_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@36445.4]
  wire  x222_inr_Foreach_sm_clock; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_reset; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_enable; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_done; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_doneLatch; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_ctrDone; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_datapathEn; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_ctrInc; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_ctrRst; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_parentAck; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_backpressure; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  x222_inr_Foreach_sm_io_break; // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36579.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36579.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36579.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36579.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36579.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@36587.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@36587.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@36587.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@36587.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@36587.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_clock; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_reset; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_wPort_0_en_0; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_full; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_active_0_in; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_active_0_out; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire [31:0] x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire [31:0] x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_rr; // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
  wire  x358_outr_UnitPipe_sm_clock; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_reset; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_enable; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_done; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_rst; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_ctrDone; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_ctrInc; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_parentAck; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  x358_outr_UnitPipe_sm_io_childAck_0; // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@36811.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@36811.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@36811.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@36811.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@36811.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@36819.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@36819.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@36819.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@36819.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@36819.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_clock; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_reset; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TVALID; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TREADY; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire [255:0] x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TDATA; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TVALID; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TREADY; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire [255:0] x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TDATA; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire [7:0] x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TID; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire [7:0] x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TDEST; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_rr; // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
  wire  _T_254; // @[package.scala 96:25:@36538.4 package.scala 96:25:@36539.4]
  wire  _T_260; // @[implicits.scala 47:10:@36542.4]
  wire  _T_261; // @[sm_x359_outr_UnitPipe.scala 70:41:@36543.4]
  wire  _T_262; // @[sm_x359_outr_UnitPipe.scala 70:78:@36544.4]
  wire  _T_263; // @[sm_x359_outr_UnitPipe.scala 70:76:@36545.4]
  wire  _T_275; // @[package.scala 96:25:@36584.4 package.scala 96:25:@36585.4]
  wire  _T_281; // @[package.scala 96:25:@36592.4 package.scala 96:25:@36593.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@36595.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@36604.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@36605.4]
  wire  _T_354; // @[package.scala 100:49:@36782.4]
  reg  _T_357; // @[package.scala 48:56:@36783.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@36816.4 package.scala 96:25:@36817.4]
  wire  _T_377; // @[package.scala 96:25:@36824.4 package.scala 96:25:@36825.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@36827.4]
  x204_fifoinraw_0 x204_fifoinraw_0 ( // @[m_x204_fifoinraw_0.scala 27:17:@36373.4]
    .clock(x204_fifoinraw_0_clock),
    .reset(x204_fifoinraw_0_reset)
  );
  x205_fifoinpacked_0 x205_fifoinpacked_0 ( // @[m_x205_fifoinpacked_0.scala 27:17:@36397.4]
    .clock(x205_fifoinpacked_0_clock),
    .reset(x205_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x205_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x205_fifoinpacked_0_io_full),
    .io_active_0_in(x205_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x205_fifoinpacked_0_io_active_0_out)
  );
  x204_fifoinraw_0 x206_fifooutraw_0 ( // @[m_x206_fifooutraw_0.scala 27:17:@36421.4]
    .clock(x206_fifooutraw_0_clock),
    .reset(x206_fifooutraw_0_reset)
  );
  x209_ctrchain x209_ctrchain ( // @[SpatialBlocks.scala 37:22:@36445.4]
    .clock(x209_ctrchain_clock),
    .reset(x209_ctrchain_reset),
    .io_input_reset(x209_ctrchain_io_input_reset),
    .io_input_enable(x209_ctrchain_io_input_enable),
    .io_output_counts_1(x209_ctrchain_io_output_counts_1),
    .io_output_counts_0(x209_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x209_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x209_ctrchain_io_output_oobs_1),
    .io_output_done(x209_ctrchain_io_output_done)
  );
  x222_inr_Foreach_sm x222_inr_Foreach_sm ( // @[sm_x222_inr_Foreach.scala 32:18:@36505.4]
    .clock(x222_inr_Foreach_sm_clock),
    .reset(x222_inr_Foreach_sm_reset),
    .io_enable(x222_inr_Foreach_sm_io_enable),
    .io_done(x222_inr_Foreach_sm_io_done),
    .io_doneLatch(x222_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x222_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x222_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x222_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x222_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x222_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x222_inr_Foreach_sm_io_backpressure),
    .io_break(x222_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36533.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36579.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@36587.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x222_inr_Foreach_kernelx222_inr_Foreach_concrete1 x222_inr_Foreach_kernelx222_inr_Foreach_concrete1 ( // @[sm_x222_inr_Foreach.scala 92:24:@36622.4]
    .clock(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_clock),
    .reset(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_reset),
    .io_in_x205_fifoinpacked_0_wPort_0_en_0(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_wPort_0_en_0),
    .io_in_x205_fifoinpacked_0_full(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_full),
    .io_in_x205_fifoinpacked_0_active_0_in(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_active_0_in),
    .io_in_x205_fifoinpacked_0_active_0_out(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x358_outr_UnitPipe_sm ( // @[sm_x358_outr_UnitPipe.scala 32:18:@36754.4]
    .clock(x358_outr_UnitPipe_sm_clock),
    .reset(x358_outr_UnitPipe_sm_reset),
    .io_enable(x358_outr_UnitPipe_sm_io_enable),
    .io_done(x358_outr_UnitPipe_sm_io_done),
    .io_rst(x358_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x358_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x358_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x358_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x358_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x358_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x358_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@36811.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@36819.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1 x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1 ( // @[sm_x358_outr_UnitPipe.scala 76:24:@36849.4]
    .clock(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_clock),
    .reset(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_reset),
    .io_in_x202_TVALID(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TVALID),
    .io_in_x202_TREADY(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TREADY),
    .io_in_x202_TDATA(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TDATA),
    .io_in_x201_TVALID(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TVALID),
    .io_in_x201_TREADY(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TREADY),
    .io_in_x201_TDATA(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TDATA),
    .io_in_x201_TID(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TID),
    .io_in_x201_TDEST(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TDEST),
    .io_sigsIn_smEnableOuts_0(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@36538.4 package.scala 96:25:@36539.4]
  assign _T_260 = x205_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@36542.4]
  assign _T_261 = ~ _T_260; // @[sm_x359_outr_UnitPipe.scala 70:41:@36543.4]
  assign _T_262 = ~ x205_fifoinpacked_0_io_active_0_out; // @[sm_x359_outr_UnitPipe.scala 70:78:@36544.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x359_outr_UnitPipe.scala 70:76:@36545.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36584.4 package.scala 96:25:@36585.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@36592.4 package.scala 96:25:@36593.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@36595.4]
  assign _T_286 = x222_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@36604.4]
  assign _T_287 = ~ x222_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@36605.4]
  assign _T_354 = x358_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@36782.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@36816.4 package.scala 96:25:@36817.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@36824.4 package.scala 96:25:@36825.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@36827.4]
  assign io_in_x202_TVALID = x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TVALID; // @[sm_x358_outr_UnitPipe.scala 48:23:@36906.4]
  assign io_in_x202_TDATA = x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TDATA; // @[sm_x358_outr_UnitPipe.scala 48:23:@36904.4]
  assign io_in_x201_TREADY = x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TREADY; // @[sm_x358_outr_UnitPipe.scala 49:23:@36914.4]
  assign io_sigsOut_smDoneIn_0 = x222_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@36602.4]
  assign io_sigsOut_smDoneIn_1 = x358_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@36834.4]
  assign io_sigsOut_smCtrCopyDone_0 = x222_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@36621.4]
  assign io_sigsOut_smCtrCopyDone_1 = x358_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@36848.4]
  assign x204_fifoinraw_0_clock = clock; // @[:@36374.4]
  assign x204_fifoinraw_0_reset = reset; // @[:@36375.4]
  assign x205_fifoinpacked_0_clock = clock; // @[:@36398.4]
  assign x205_fifoinpacked_0_reset = reset; // @[:@36399.4]
  assign x205_fifoinpacked_0_io_wPort_0_en_0 = x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@36682.4]
  assign x205_fifoinpacked_0_io_active_0_in = x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@36681.4]
  assign x206_fifooutraw_0_clock = clock; // @[:@36422.4]
  assign x206_fifooutraw_0_reset = reset; // @[:@36423.4]
  assign x209_ctrchain_clock = clock; // @[:@36446.4]
  assign x209_ctrchain_reset = reset; // @[:@36447.4]
  assign x209_ctrchain_io_input_reset = x222_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@36620.4]
  assign x209_ctrchain_io_input_enable = x222_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@36572.4 SpatialBlocks.scala 159:42:@36619.4]
  assign x222_inr_Foreach_sm_clock = clock; // @[:@36506.4]
  assign x222_inr_Foreach_sm_reset = reset; // @[:@36507.4]
  assign x222_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@36599.4]
  assign x222_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x359_outr_UnitPipe.scala 69:38:@36541.4]
  assign x222_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@36601.4]
  assign x222_inr_Foreach_sm_io_backpressure = _T_263 | x222_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@36573.4]
  assign x222_inr_Foreach_sm_io_break = 1'h0; // @[sm_x359_outr_UnitPipe.scala 73:36:@36551.4]
  assign RetimeWrapper_clock = clock; // @[:@36534.4]
  assign RetimeWrapper_reset = reset; // @[:@36535.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36537.4]
  assign RetimeWrapper_io_in = x209_ctrchain_io_output_done; // @[package.scala 94:16:@36536.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36580.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36581.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36583.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@36582.4]
  assign RetimeWrapper_2_clock = clock; // @[:@36588.4]
  assign RetimeWrapper_2_reset = reset; // @[:@36589.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@36591.4]
  assign RetimeWrapper_2_io_in = x222_inr_Foreach_sm_io_done; // @[package.scala 94:16:@36590.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_clock = clock; // @[:@36623.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_reset = reset; // @[:@36624.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_full = x205_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@36676.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_in_x205_fifoinpacked_0_active_0_out = x205_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@36675.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x222_inr_Foreach_sm_io_doneLatch; // @[sm_x222_inr_Foreach.scala 97:22:@36705.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x222_inr_Foreach.scala 97:22:@36703.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_break = x222_inr_Foreach_sm_io_break; // @[sm_x222_inr_Foreach.scala 97:22:@36701.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x209_ctrchain_io_output_counts_1[12]}},x209_ctrchain_io_output_counts_1}; // @[sm_x222_inr_Foreach.scala 97:22:@36696.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x209_ctrchain_io_output_counts_0[12]}},x209_ctrchain_io_output_counts_0}; // @[sm_x222_inr_Foreach.scala 97:22:@36695.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x209_ctrchain_io_output_oobs_0; // @[sm_x222_inr_Foreach.scala 97:22:@36693.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x209_ctrchain_io_output_oobs_1; // @[sm_x222_inr_Foreach.scala 97:22:@36694.4]
  assign x222_inr_Foreach_kernelx222_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x222_inr_Foreach.scala 96:18:@36689.4]
  assign x358_outr_UnitPipe_sm_clock = clock; // @[:@36755.4]
  assign x358_outr_UnitPipe_sm_reset = reset; // @[:@36756.4]
  assign x358_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@36831.4]
  assign x358_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@36806.4]
  assign x358_outr_UnitPipe_sm_io_ctrDone = x358_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x359_outr_UnitPipe.scala 78:40:@36786.4]
  assign x358_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@36833.4]
  assign x358_outr_UnitPipe_sm_io_doneIn_0 = x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@36803.4]
  assign RetimeWrapper_3_clock = clock; // @[:@36812.4]
  assign RetimeWrapper_3_reset = reset; // @[:@36813.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@36815.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@36814.4]
  assign RetimeWrapper_4_clock = clock; // @[:@36820.4]
  assign RetimeWrapper_4_reset = reset; // @[:@36821.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@36823.4]
  assign RetimeWrapper_4_io_in = x358_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@36822.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_clock = clock; // @[:@36850.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_reset = reset; // @[:@36851.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x202_TREADY = io_in_x202_TREADY; // @[sm_x358_outr_UnitPipe.scala 48:23:@36905.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TVALID = io_in_x201_TVALID; // @[sm_x358_outr_UnitPipe.scala 49:23:@36915.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TDATA = io_in_x201_TDATA; // @[sm_x358_outr_UnitPipe.scala 49:23:@36913.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TID = io_in_x201_TID; // @[sm_x358_outr_UnitPipe.scala 49:23:@36909.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_in_x201_TDEST = io_in_x201_TDEST; // @[sm_x358_outr_UnitPipe.scala 49:23:@36908.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x358_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x358_outr_UnitPipe.scala 81:22:@36924.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x358_outr_UnitPipe_sm_io_childAck_0; // @[sm_x358_outr_UnitPipe.scala 81:22:@36922.4]
  assign x358_outr_UnitPipe_kernelx358_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x358_outr_UnitPipe.scala 80:18:@36916.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x381_outr_UnitPipe_sm( // @[:@37413.2]
  input   clock, // @[:@37414.4]
  input   reset, // @[:@37415.4]
  input   io_enable, // @[:@37416.4]
  output  io_done, // @[:@37416.4]
  input   io_parentAck, // @[:@37416.4]
  input   io_doneIn_0, // @[:@37416.4]
  input   io_doneIn_1, // @[:@37416.4]
  input   io_doneIn_2, // @[:@37416.4]
  output  io_enableOut_0, // @[:@37416.4]
  output  io_enableOut_1, // @[:@37416.4]
  output  io_enableOut_2, // @[:@37416.4]
  output  io_childAck_0, // @[:@37416.4]
  output  io_childAck_1, // @[:@37416.4]
  output  io_childAck_2, // @[:@37416.4]
  input   io_ctrCopyDone_0, // @[:@37416.4]
  input   io_ctrCopyDone_1, // @[:@37416.4]
  input   io_ctrCopyDone_2 // @[:@37416.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@37419.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@37419.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@37419.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@37419.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@37419.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@37419.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@37422.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@37422.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@37422.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@37422.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@37422.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@37422.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@37425.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@37425.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@37425.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@37425.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@37425.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@37425.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@37428.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@37428.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@37428.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@37428.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@37428.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@37428.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@37431.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@37431.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@37431.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@37431.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@37431.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@37431.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@37434.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@37434.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@37434.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@37434.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@37434.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@37434.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@37475.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@37475.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@37475.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@37475.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@37475.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@37475.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@37478.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@37478.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@37478.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@37478.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@37478.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@37478.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@37481.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@37481.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@37481.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@37481.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@37481.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@37481.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37532.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37532.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37532.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37532.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37532.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37546.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37546.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37546.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37546.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37546.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@37564.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@37564.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@37564.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@37564.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@37564.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@37615.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@37615.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@37615.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@37615.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@37615.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@37633.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@37633.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@37633.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@37633.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@37633.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@37684.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@37684.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@37684.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@37684.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@37684.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@37702.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@37702.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@37702.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@37702.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@37702.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@37759.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@37759.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@37759.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@37759.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@37759.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@37776.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@37776.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@37776.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@37776.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@37776.4]
  wire  _T_77; // @[Controllers.scala 80:47:@37437.4]
  wire  allDone; // @[Controllers.scala 80:47:@37438.4]
  wire  _T_151; // @[Controllers.scala 165:35:@37516.4]
  wire  _T_153; // @[Controllers.scala 165:60:@37517.4]
  wire  _T_154; // @[Controllers.scala 165:58:@37518.4]
  wire  _T_156; // @[Controllers.scala 165:76:@37519.4]
  wire  _T_157; // @[Controllers.scala 165:74:@37520.4]
  wire  _T_161; // @[Controllers.scala 165:109:@37523.4]
  wire  _T_164; // @[Controllers.scala 165:141:@37525.4]
  wire  _T_172; // @[package.scala 96:25:@37537.4 package.scala 96:25:@37538.4]
  wire  _T_176; // @[Controllers.scala 167:54:@37540.4]
  wire  _T_177; // @[Controllers.scala 167:52:@37541.4]
  wire  _T_184; // @[package.scala 96:25:@37551.4 package.scala 96:25:@37552.4]
  wire  _T_202; // @[package.scala 96:25:@37569.4 package.scala 96:25:@37570.4]
  wire  _T_206; // @[Controllers.scala 169:67:@37572.4]
  wire  _T_207; // @[Controllers.scala 169:86:@37573.4]
  wire  _T_219; // @[Controllers.scala 165:35:@37585.4]
  wire  _T_221; // @[Controllers.scala 165:60:@37586.4]
  wire  _T_222; // @[Controllers.scala 165:58:@37587.4]
  wire  _T_224; // @[Controllers.scala 165:76:@37588.4]
  wire  _T_225; // @[Controllers.scala 165:74:@37589.4]
  wire  _T_229; // @[Controllers.scala 165:109:@37592.4]
  wire  _T_232; // @[Controllers.scala 165:141:@37594.4]
  wire  _T_240; // @[package.scala 96:25:@37606.4 package.scala 96:25:@37607.4]
  wire  _T_244; // @[Controllers.scala 167:54:@37609.4]
  wire  _T_245; // @[Controllers.scala 167:52:@37610.4]
  wire  _T_252; // @[package.scala 96:25:@37620.4 package.scala 96:25:@37621.4]
  wire  _T_270; // @[package.scala 96:25:@37638.4 package.scala 96:25:@37639.4]
  wire  _T_274; // @[Controllers.scala 169:67:@37641.4]
  wire  _T_275; // @[Controllers.scala 169:86:@37642.4]
  wire  _T_287; // @[Controllers.scala 165:35:@37654.4]
  wire  _T_289; // @[Controllers.scala 165:60:@37655.4]
  wire  _T_290; // @[Controllers.scala 165:58:@37656.4]
  wire  _T_292; // @[Controllers.scala 165:76:@37657.4]
  wire  _T_293; // @[Controllers.scala 165:74:@37658.4]
  wire  _T_297; // @[Controllers.scala 165:109:@37661.4]
  wire  _T_300; // @[Controllers.scala 165:141:@37663.4]
  wire  _T_308; // @[package.scala 96:25:@37675.4 package.scala 96:25:@37676.4]
  wire  _T_312; // @[Controllers.scala 167:54:@37678.4]
  wire  _T_313; // @[Controllers.scala 167:52:@37679.4]
  wire  _T_320; // @[package.scala 96:25:@37689.4 package.scala 96:25:@37690.4]
  wire  _T_338; // @[package.scala 96:25:@37707.4 package.scala 96:25:@37708.4]
  wire  _T_342; // @[Controllers.scala 169:67:@37710.4]
  wire  _T_343; // @[Controllers.scala 169:86:@37711.4]
  wire  _T_358; // @[Controllers.scala 213:68:@37729.4]
  wire  _T_360; // @[Controllers.scala 213:90:@37731.4]
  wire  _T_362; // @[Controllers.scala 213:132:@37733.4]
  wire  _T_366; // @[Controllers.scala 213:68:@37738.4]
  wire  _T_368; // @[Controllers.scala 213:90:@37740.4]
  wire  _T_374; // @[Controllers.scala 213:68:@37746.4]
  wire  _T_376; // @[Controllers.scala 213:90:@37748.4]
  wire  _T_383; // @[package.scala 100:49:@37754.4]
  reg  _T_386; // @[package.scala 48:56:@37755.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@37757.4]
  reg  _T_400; // @[package.scala 48:56:@37773.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@37419.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@37422.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@37425.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@37428.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@37431.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@37434.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@37475.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@37478.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@37481.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@37532.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@37546.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@37564.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@37601.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@37615.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@37633.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@37670.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@37684.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@37702.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@37759.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@37776.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@37437.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@37438.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@37516.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@37517.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@37518.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@37519.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@37520.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@37523.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@37525.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@37537.4 package.scala 96:25:@37538.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@37540.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@37541.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37551.4 package.scala 96:25:@37552.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@37569.4 package.scala 96:25:@37570.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@37572.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@37573.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@37585.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@37586.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@37587.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@37588.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@37589.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@37592.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@37594.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@37606.4 package.scala 96:25:@37607.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@37609.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@37610.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@37620.4 package.scala 96:25:@37621.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@37638.4 package.scala 96:25:@37639.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@37641.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@37642.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@37654.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@37655.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@37656.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@37657.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@37658.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@37661.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@37663.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@37675.4 package.scala 96:25:@37676.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@37678.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@37679.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@37689.4 package.scala 96:25:@37690.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@37707.4 package.scala 96:25:@37708.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@37710.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@37711.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@37729.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@37731.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@37733.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@37738.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@37740.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@37746.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@37748.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@37754.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@37757.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@37783.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@37737.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@37745.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@37753.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@37724.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@37726.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@37728.4]
  assign active_0_clock = clock; // @[:@37420.4]
  assign active_0_reset = reset; // @[:@37421.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@37527.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@37531.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@37441.4]
  assign active_1_clock = clock; // @[:@37423.4]
  assign active_1_reset = reset; // @[:@37424.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@37596.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@37600.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@37442.4]
  assign active_2_clock = clock; // @[:@37426.4]
  assign active_2_reset = reset; // @[:@37427.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@37665.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@37669.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@37443.4]
  assign done_0_clock = clock; // @[:@37429.4]
  assign done_0_reset = reset; // @[:@37430.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@37577.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@37455.4 Controllers.scala 170:32:@37584.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@37444.4]
  assign done_1_clock = clock; // @[:@37432.4]
  assign done_1_reset = reset; // @[:@37433.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@37646.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@37464.4 Controllers.scala 170:32:@37653.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@37445.4]
  assign done_2_clock = clock; // @[:@37435.4]
  assign done_2_reset = reset; // @[:@37436.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@37715.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@37473.4 Controllers.scala 170:32:@37722.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@37446.4]
  assign iterDone_0_clock = clock; // @[:@37476.4]
  assign iterDone_0_reset = reset; // @[:@37477.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@37545.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@37495.4 Controllers.scala 168:36:@37561.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@37484.4]
  assign iterDone_1_clock = clock; // @[:@37479.4]
  assign iterDone_1_reset = reset; // @[:@37480.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@37614.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@37504.4 Controllers.scala 168:36:@37630.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@37485.4]
  assign iterDone_2_clock = clock; // @[:@37482.4]
  assign iterDone_2_reset = reset; // @[:@37483.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@37683.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@37513.4 Controllers.scala 168:36:@37699.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@37486.4]
  assign RetimeWrapper_clock = clock; // @[:@37533.4]
  assign RetimeWrapper_reset = reset; // @[:@37534.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@37536.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@37535.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37547.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37548.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@37550.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@37549.4]
  assign RetimeWrapper_2_clock = clock; // @[:@37565.4]
  assign RetimeWrapper_2_reset = reset; // @[:@37566.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@37568.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@37567.4]
  assign RetimeWrapper_3_clock = clock; // @[:@37602.4]
  assign RetimeWrapper_3_reset = reset; // @[:@37603.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@37605.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@37604.4]
  assign RetimeWrapper_4_clock = clock; // @[:@37616.4]
  assign RetimeWrapper_4_reset = reset; // @[:@37617.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@37619.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@37618.4]
  assign RetimeWrapper_5_clock = clock; // @[:@37634.4]
  assign RetimeWrapper_5_reset = reset; // @[:@37635.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@37637.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@37636.4]
  assign RetimeWrapper_6_clock = clock; // @[:@37671.4]
  assign RetimeWrapper_6_reset = reset; // @[:@37672.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@37674.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@37673.4]
  assign RetimeWrapper_7_clock = clock; // @[:@37685.4]
  assign RetimeWrapper_7_reset = reset; // @[:@37686.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@37688.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@37687.4]
  assign RetimeWrapper_8_clock = clock; // @[:@37703.4]
  assign RetimeWrapper_8_reset = reset; // @[:@37704.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@37706.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@37705.4]
  assign RetimeWrapper_9_clock = clock; // @[:@37760.4]
  assign RetimeWrapper_9_reset = reset; // @[:@37761.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@37763.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@37762.4]
  assign RetimeWrapper_10_clock = clock; // @[:@37777.4]
  assign RetimeWrapper_10_reset = reset; // @[:@37778.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@37780.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@37779.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x367_inr_UnitPipe_sm( // @[:@37956.2]
  input   clock, // @[:@37957.4]
  input   reset, // @[:@37958.4]
  input   io_enable, // @[:@37959.4]
  output  io_done, // @[:@37959.4]
  output  io_doneLatch, // @[:@37959.4]
  input   io_ctrDone, // @[:@37959.4]
  output  io_datapathEn, // @[:@37959.4]
  output  io_ctrInc, // @[:@37959.4]
  input   io_parentAck, // @[:@37959.4]
  input   io_backpressure // @[:@37959.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@37961.4]
  wire  active_reset; // @[Controllers.scala 261:22:@37961.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@37961.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@37961.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@37961.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@37961.4]
  wire  done_clock; // @[Controllers.scala 262:20:@37964.4]
  wire  done_reset; // @[Controllers.scala 262:20:@37964.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@37964.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@37964.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@37964.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@37964.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38018.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38018.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38018.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38018.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38018.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38026.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38026.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38026.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38026.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38026.4]
  wire  _T_80; // @[Controllers.scala 264:48:@37969.4]
  wire  _T_81; // @[Controllers.scala 264:46:@37970.4]
  wire  _T_82; // @[Controllers.scala 264:62:@37971.4]
  wire  _T_83; // @[Controllers.scala 264:60:@37972.4]
  wire  _T_100; // @[package.scala 100:49:@37989.4]
  reg  _T_103; // @[package.scala 48:56:@37990.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@37998.4]
  wire  _T_116; // @[Controllers.scala 283:41:@38006.4]
  wire  _T_117; // @[Controllers.scala 283:59:@38007.4]
  wire  _T_119; // @[Controllers.scala 284:37:@38010.4]
  reg  _T_125; // @[package.scala 48:56:@38014.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@38036.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@38039.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@38041.4]
  wire  _T_152; // @[Controllers.scala 292:61:@38042.4]
  wire  _T_153; // @[Controllers.scala 292:24:@38043.4]
  SRFF active ( // @[Controllers.scala 261:22:@37961.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@37964.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@38018.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@38026.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@37969.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@37970.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@37971.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@37972.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@37989.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@37998.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@38006.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@38007.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@38010.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@38041.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@38042.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@38043.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@38017.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@38045.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@38009.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@38012.4]
  assign active_clock = clock; // @[:@37962.4]
  assign active_reset = reset; // @[:@37963.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@37974.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@37978.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@37979.4]
  assign done_clock = clock; // @[:@37965.4]
  assign done_reset = reset; // @[:@37966.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@37994.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@37987.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@37988.4]
  assign RetimeWrapper_clock = clock; // @[:@38019.4]
  assign RetimeWrapper_reset = reset; // @[:@38020.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@38022.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@38021.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38027.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38028.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@38030.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@38029.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1( // @[:@38120.2]
  output        io_in_x360_valid, // @[:@38123.4]
  output [63:0] io_in_x360_bits_addr, // @[:@38123.4]
  output [31:0] io_in_x360_bits_size, // @[:@38123.4]
  input  [63:0] io_in_x199_outdram_number, // @[:@38123.4]
  input         io_sigsIn_backpressure, // @[:@38123.4]
  input         io_sigsIn_datapathEn, // @[:@38123.4]
  input         io_rr // @[:@38123.4]
);
  wire [96:0] x364_tuple; // @[Cat.scala 30:58:@38137.4]
  wire  _T_135; // @[implicits.scala 55:10:@38140.4]
  assign x364_tuple = {33'h7e9000,io_in_x199_outdram_number}; // @[Cat.scala 30:58:@38137.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@38140.4]
  assign io_in_x360_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x367_inr_UnitPipe.scala 65:18:@38143.4]
  assign io_in_x360_bits_addr = x364_tuple[63:0]; // @[sm_x367_inr_UnitPipe.scala 66:22:@38145.4]
  assign io_in_x360_bits_size = x364_tuple[95:64]; // @[sm_x367_inr_UnitPipe.scala 67:22:@38147.4]
endmodule
module FF_13( // @[:@38149.2]
  input         clock, // @[:@38150.4]
  input         reset, // @[:@38151.4]
  output [22:0] io_rPort_0_output_0, // @[:@38152.4]
  input  [22:0] io_wPort_0_data_0, // @[:@38152.4]
  input         io_wPort_0_reset, // @[:@38152.4]
  input         io_wPort_0_en_0 // @[:@38152.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@38167.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@38169.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@38170.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@38169.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@38170.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@38172.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@38187.2]
  input         clock, // @[:@38188.4]
  input         reset, // @[:@38189.4]
  input         io_input_reset, // @[:@38190.4]
  input         io_input_enable, // @[:@38190.4]
  output [22:0] io_output_count_0, // @[:@38190.4]
  output        io_output_oobs_0, // @[:@38190.4]
  output        io_output_done // @[:@38190.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@38203.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@38203.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@38203.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@38203.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@38203.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@38203.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@38219.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@38219.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@38219.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@38219.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@38219.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@38219.4]
  wire  _T_36; // @[Counter.scala 264:45:@38222.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@38247.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@38248.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@38249.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@38250.4]
  wire  _T_57; // @[Counter.scala 293:18:@38252.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@38260.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@38263.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@38264.4]
  wire  _T_75; // @[Counter.scala 322:102:@38268.4]
  wire  _T_77; // @[Counter.scala 322:130:@38269.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@38203.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@38219.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@38222.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@38247.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@38248.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@38249.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@38250.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@38252.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@38260.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@38263.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@38264.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@38268.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@38269.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@38267.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@38271.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@38273.4]
  assign bases_0_clock = clock; // @[:@38204.4]
  assign bases_0_reset = reset; // @[:@38205.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@38266.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@38245.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@38246.4]
  assign SRFF_clock = clock; // @[:@38220.4]
  assign SRFF_reset = reset; // @[:@38221.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@38224.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@38226.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@38227.4]
endmodule
module x369_ctrchain( // @[:@38278.2]
  input         clock, // @[:@38279.4]
  input         reset, // @[:@38280.4]
  input         io_input_reset, // @[:@38281.4]
  input         io_input_enable, // @[:@38281.4]
  output [22:0] io_output_counts_0, // @[:@38281.4]
  output        io_output_oobs_0, // @[:@38281.4]
  output        io_output_done // @[:@38281.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@38283.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@38283.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@38283.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@38283.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@38283.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@38283.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@38283.4]
  reg  wasDone; // @[Counter.scala 542:24:@38292.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@38298.4]
  wire  _T_47; // @[Counter.scala 546:80:@38299.4]
  reg  doneLatch; // @[Counter.scala 550:26:@38304.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@38305.4]
  wire  _T_55; // @[Counter.scala 551:19:@38306.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@38283.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@38298.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@38299.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@38305.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@38306.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@38308.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@38310.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@38301.4]
  assign ctrs_0_clock = clock; // @[:@38284.4]
  assign ctrs_0_reset = reset; // @[:@38285.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@38289.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@38290.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x376_inr_Foreach_sm( // @[:@38498.2]
  input   clock, // @[:@38499.4]
  input   reset, // @[:@38500.4]
  input   io_enable, // @[:@38501.4]
  output  io_done, // @[:@38501.4]
  output  io_doneLatch, // @[:@38501.4]
  input   io_ctrDone, // @[:@38501.4]
  output  io_datapathEn, // @[:@38501.4]
  output  io_ctrInc, // @[:@38501.4]
  output  io_ctrRst, // @[:@38501.4]
  input   io_parentAck, // @[:@38501.4]
  input   io_backpressure, // @[:@38501.4]
  input   io_break // @[:@38501.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@38503.4]
  wire  active_reset; // @[Controllers.scala 261:22:@38503.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@38503.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@38503.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@38503.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@38503.4]
  wire  done_clock; // @[Controllers.scala 262:20:@38506.4]
  wire  done_reset; // @[Controllers.scala 262:20:@38506.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@38506.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@38506.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@38506.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@38506.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38540.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38540.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38540.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38540.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38540.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38562.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38562.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38562.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38562.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38562.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38574.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38574.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38574.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@38574.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@38574.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38582.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38582.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38582.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@38582.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@38582.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@38598.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@38598.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@38598.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@38598.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@38598.4]
  wire  _T_80; // @[Controllers.scala 264:48:@38511.4]
  wire  _T_81; // @[Controllers.scala 264:46:@38512.4]
  wire  _T_82; // @[Controllers.scala 264:62:@38513.4]
  wire  _T_83; // @[Controllers.scala 264:60:@38514.4]
  wire  _T_100; // @[package.scala 100:49:@38531.4]
  reg  _T_103; // @[package.scala 48:56:@38532.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@38545.4 package.scala 96:25:@38546.4]
  wire  _T_110; // @[package.scala 100:49:@38547.4]
  reg  _T_113; // @[package.scala 48:56:@38548.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@38550.4]
  wire  _T_118; // @[Controllers.scala 283:41:@38555.4]
  wire  _T_119; // @[Controllers.scala 283:59:@38556.4]
  wire  _T_121; // @[Controllers.scala 284:37:@38559.4]
  wire  _T_124; // @[package.scala 96:25:@38567.4 package.scala 96:25:@38568.4]
  wire  _T_126; // @[package.scala 100:49:@38569.4]
  reg  _T_129; // @[package.scala 48:56:@38570.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@38592.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@38594.4]
  reg  _T_153; // @[package.scala 48:56:@38595.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@38603.4 package.scala 96:25:@38604.4]
  wire  _T_158; // @[Controllers.scala 292:61:@38605.4]
  wire  _T_159; // @[Controllers.scala 292:24:@38606.4]
  SRFF active ( // @[Controllers.scala 261:22:@38503.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@38506.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@38540.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@38562.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@38574.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@38582.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@38598.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@38511.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@38512.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@38513.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@38514.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@38531.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@38545.4 package.scala 96:25:@38546.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@38547.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@38550.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@38555.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@38556.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@38559.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@38567.4 package.scala 96:25:@38568.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@38569.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@38594.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@38603.4 package.scala 96:25:@38604.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@38605.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@38606.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@38573.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@38608.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@38558.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@38561.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@38553.4]
  assign active_clock = clock; // @[:@38504.4]
  assign active_reset = reset; // @[:@38505.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@38516.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@38520.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@38521.4]
  assign done_clock = clock; // @[:@38507.4]
  assign done_reset = reset; // @[:@38508.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@38536.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@38529.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@38530.4]
  assign RetimeWrapper_clock = clock; // @[:@38541.4]
  assign RetimeWrapper_reset = reset; // @[:@38542.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@38544.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@38543.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38563.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38564.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@38566.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@38565.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38575.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38576.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@38578.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@38577.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38583.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38584.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@38586.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@38585.4]
  assign RetimeWrapper_4_clock = clock; // @[:@38599.4]
  assign RetimeWrapper_4_reset = reset; // @[:@38600.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@38602.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@38601.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x376_inr_Foreach_kernelx376_inr_Foreach_concrete1( // @[:@38815.2]
  input         clock, // @[:@38816.4]
  input         reset, // @[:@38817.4]
  output        io_in_x361_valid, // @[:@38818.4]
  output [31:0] io_in_x361_bits_wdata_0, // @[:@38818.4]
  output        io_in_x361_bits_wstrb, // @[:@38818.4]
  output [20:0] io_in_x203_outbuf_0_rPort_0_ofs_0, // @[:@38818.4]
  output        io_in_x203_outbuf_0_rPort_0_en_0, // @[:@38818.4]
  output        io_in_x203_outbuf_0_rPort_0_backpressure, // @[:@38818.4]
  input  [31:0] io_in_x203_outbuf_0_rPort_0_output_0, // @[:@38818.4]
  input         io_sigsIn_backpressure, // @[:@38818.4]
  input         io_sigsIn_datapathEn, // @[:@38818.4]
  input         io_sigsIn_break, // @[:@38818.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@38818.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@38818.4]
  input         io_rr // @[:@38818.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@38845.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@38845.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38874.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38874.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38874.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38874.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38874.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38883.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38883.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38883.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38883.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38883.4]
  wire  b371; // @[sm_x376_inr_Foreach.scala 62:18:@38853.4]
  wire  _T_274; // @[sm_x376_inr_Foreach.scala 67:129:@38857.4]
  wire  _T_278; // @[implicits.scala 55:10:@38860.4]
  wire  _T_279; // @[sm_x376_inr_Foreach.scala 67:146:@38861.4]
  wire [32:0] x374_tuple; // @[Cat.scala 30:58:@38871.4]
  wire  _T_290; // @[package.scala 96:25:@38888.4 package.scala 96:25:@38889.4]
  wire  _T_292; // @[implicits.scala 55:10:@38890.4]
  wire  x561_b371_D2; // @[package.scala 96:25:@38879.4 package.scala 96:25:@38880.4]
  wire  _T_293; // @[sm_x376_inr_Foreach.scala 74:112:@38891.4]
  wire [31:0] b370_number; // @[Math.scala 723:22:@38850.4 Math.scala 724:14:@38851.4]
  _ _ ( // @[Math.scala 720:24:@38845.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@38874.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@38883.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b371 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x376_inr_Foreach.scala 62:18:@38853.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x376_inr_Foreach.scala 67:129:@38857.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@38860.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x376_inr_Foreach.scala 67:146:@38861.4]
  assign x374_tuple = {1'h1,io_in_x203_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@38871.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@38888.4 package.scala 96:25:@38889.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@38890.4]
  assign x561_b371_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@38879.4 package.scala 96:25:@38880.4]
  assign _T_293 = _T_292 & x561_b371_D2; // @[sm_x376_inr_Foreach.scala 74:112:@38891.4]
  assign b370_number = __io_result; // @[Math.scala 723:22:@38850.4 Math.scala 724:14:@38851.4]
  assign io_in_x361_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x376_inr_Foreach.scala 74:18:@38893.4]
  assign io_in_x361_bits_wdata_0 = x374_tuple[31:0]; // @[sm_x376_inr_Foreach.scala 75:26:@38895.4]
  assign io_in_x361_bits_wstrb = x374_tuple[32]; // @[sm_x376_inr_Foreach.scala 76:23:@38897.4]
  assign io_in_x203_outbuf_0_rPort_0_ofs_0 = b370_number[20:0]; // @[MemInterfaceType.scala 107:54:@38864.4]
  assign io_in_x203_outbuf_0_rPort_0_en_0 = _T_279 & b371; // @[MemInterfaceType.scala 110:79:@38866.4]
  assign io_in_x203_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38865.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@38848.4]
  assign RetimeWrapper_clock = clock; // @[:@38875.4]
  assign RetimeWrapper_reset = reset; // @[:@38876.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38878.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@38877.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38884.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38885.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38887.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38886.4]
endmodule
module x380_inr_UnitPipe_sm( // @[:@39053.2]
  input   clock, // @[:@39054.4]
  input   reset, // @[:@39055.4]
  input   io_enable, // @[:@39056.4]
  output  io_done, // @[:@39056.4]
  output  io_doneLatch, // @[:@39056.4]
  input   io_ctrDone, // @[:@39056.4]
  output  io_datapathEn, // @[:@39056.4]
  output  io_ctrInc, // @[:@39056.4]
  input   io_parentAck // @[:@39056.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@39058.4]
  wire  active_reset; // @[Controllers.scala 261:22:@39058.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@39058.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@39058.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@39058.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@39058.4]
  wire  done_clock; // @[Controllers.scala 262:20:@39061.4]
  wire  done_reset; // @[Controllers.scala 262:20:@39061.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@39061.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@39061.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@39061.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@39061.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39095.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39095.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39095.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39095.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39095.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39117.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39117.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39117.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39117.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39117.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@39129.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@39129.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@39129.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@39129.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@39129.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@39137.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@39137.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@39137.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@39137.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@39137.4]
  wire  _T_80; // @[Controllers.scala 264:48:@39066.4]
  wire  _T_81; // @[Controllers.scala 264:46:@39067.4]
  wire  _T_82; // @[Controllers.scala 264:62:@39068.4]
  wire  _T_100; // @[package.scala 100:49:@39086.4]
  reg  _T_103; // @[package.scala 48:56:@39087.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@39110.4]
  wire  _T_124; // @[package.scala 96:25:@39122.4 package.scala 96:25:@39123.4]
  wire  _T_126; // @[package.scala 100:49:@39124.4]
  reg  _T_129; // @[package.scala 48:56:@39125.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@39147.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@39149.4]
  reg  _T_153; // @[package.scala 48:56:@39150.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@39152.4]
  wire  _T_156; // @[Controllers.scala 292:61:@39153.4]
  wire  _T_157; // @[Controllers.scala 292:24:@39154.4]
  SRFF active ( // @[Controllers.scala 261:22:@39058.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@39061.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39095.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39117.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@39129.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@39137.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@39066.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@39067.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@39068.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@39086.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@39110.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@39122.4 package.scala 96:25:@39123.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@39124.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@39149.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@39152.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@39153.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@39154.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@39128.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@39156.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@39113.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@39116.4]
  assign active_clock = clock; // @[:@39059.4]
  assign active_reset = reset; // @[:@39060.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@39071.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@39075.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@39076.4]
  assign done_clock = clock; // @[:@39062.4]
  assign done_reset = reset; // @[:@39063.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@39091.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@39084.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@39085.4]
  assign RetimeWrapper_clock = clock; // @[:@39096.4]
  assign RetimeWrapper_reset = reset; // @[:@39097.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39099.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@39098.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39118.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39119.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39121.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@39120.4]
  assign RetimeWrapper_2_clock = clock; // @[:@39130.4]
  assign RetimeWrapper_2_reset = reset; // @[:@39131.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@39133.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@39132.4]
  assign RetimeWrapper_3_clock = clock; // @[:@39138.4]
  assign RetimeWrapper_3_reset = reset; // @[:@39139.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@39141.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@39140.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1( // @[:@39231.2]
  output  io_in_x362_ready, // @[:@39234.4]
  input   io_sigsIn_datapathEn // @[:@39234.4]
);
  assign io_in_x362_ready = io_sigsIn_datapathEn; // @[sm_x380_inr_UnitPipe.scala 57:18:@39246.4]
endmodule
module x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1( // @[:@39249.2]
  input         clock, // @[:@39250.4]
  input         reset, // @[:@39251.4]
  input         io_in_x361_ready, // @[:@39252.4]
  output        io_in_x361_valid, // @[:@39252.4]
  output [31:0] io_in_x361_bits_wdata_0, // @[:@39252.4]
  output        io_in_x361_bits_wstrb, // @[:@39252.4]
  input         io_in_x360_ready, // @[:@39252.4]
  output        io_in_x360_valid, // @[:@39252.4]
  output [63:0] io_in_x360_bits_addr, // @[:@39252.4]
  output [31:0] io_in_x360_bits_size, // @[:@39252.4]
  output        io_in_x362_ready, // @[:@39252.4]
  input         io_in_x362_valid, // @[:@39252.4]
  input  [63:0] io_in_x199_outdram_number, // @[:@39252.4]
  output [20:0] io_in_x203_outbuf_0_rPort_0_ofs_0, // @[:@39252.4]
  output        io_in_x203_outbuf_0_rPort_0_en_0, // @[:@39252.4]
  output        io_in_x203_outbuf_0_rPort_0_backpressure, // @[:@39252.4]
  input  [31:0] io_in_x203_outbuf_0_rPort_0_output_0, // @[:@39252.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@39252.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@39252.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@39252.4]
  input         io_sigsIn_smChildAcks_0, // @[:@39252.4]
  input         io_sigsIn_smChildAcks_1, // @[:@39252.4]
  input         io_sigsIn_smChildAcks_2, // @[:@39252.4]
  output        io_sigsOut_smDoneIn_0, // @[:@39252.4]
  output        io_sigsOut_smDoneIn_1, // @[:@39252.4]
  output        io_sigsOut_smDoneIn_2, // @[:@39252.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@39252.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@39252.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@39252.4]
  input         io_rr // @[:@39252.4]
);
  wire  x367_inr_UnitPipe_sm_clock; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_reset; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_enable; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_done; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_doneLatch; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_ctrDone; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_datapathEn; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_ctrInc; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_parentAck; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  x367_inr_UnitPipe_sm_io_backpressure; // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39376.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39376.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39376.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39376.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39376.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39384.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39384.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39384.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39384.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39384.4]
  wire  x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_valid; // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
  wire [63:0] x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_bits_addr; // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
  wire [31:0] x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_bits_size; // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
  wire [63:0] x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x199_outdram_number; // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
  wire  x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
  wire  x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
  wire  x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_rr; // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
  wire  x369_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@39482.4]
  wire  x369_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@39482.4]
  wire  x369_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@39482.4]
  wire  x369_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@39482.4]
  wire [22:0] x369_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@39482.4]
  wire  x369_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@39482.4]
  wire  x369_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@39482.4]
  wire  x376_inr_Foreach_sm_clock; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_reset; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_enable; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_done; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_doneLatch; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_ctrDone; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_datapathEn; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_ctrInc; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_ctrRst; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_parentAck; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_backpressure; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  x376_inr_Foreach_sm_io_break; // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@39603.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@39603.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@39603.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@39603.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@39603.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@39611.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@39611.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@39611.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@39611.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@39611.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_clock; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_reset; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_valid; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire [31:0] x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_bits_wdata_0; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_bits_wstrb; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire [20:0] x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_en_0; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire [31:0] x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_output_0; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire [31:0] x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_rr; // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
  wire  x380_inr_UnitPipe_sm_clock; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_reset; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_io_enable; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_io_done; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_io_doneLatch; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_io_ctrDone; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_io_datapathEn; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_io_ctrInc; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  x380_inr_UnitPipe_sm_io_parentAck; // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@39823.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@39823.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@39823.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@39823.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@39823.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@39831.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@39831.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@39831.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@39831.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@39831.4]
  wire  x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1_io_in_x362_ready; // @[sm_x380_inr_UnitPipe.scala 60:24:@39861.4]
  wire  x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x380_inr_UnitPipe.scala 60:24:@39861.4]
  wire  _T_359; // @[package.scala 100:49:@39347.4]
  reg  _T_362; // @[package.scala 48:56:@39348.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@39381.4 package.scala 96:25:@39382.4]
  wire  _T_381; // @[package.scala 96:25:@39389.4 package.scala 96:25:@39390.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@39392.4]
  wire  _T_454; // @[package.scala 96:25:@39568.4 package.scala 96:25:@39569.4]
  wire  _T_468; // @[package.scala 96:25:@39608.4 package.scala 96:25:@39609.4]
  wire  _T_474; // @[package.scala 96:25:@39616.4 package.scala 96:25:@39617.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@39619.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@39628.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@39629.4]
  wire  _T_547; // @[package.scala 100:49:@39794.4]
  reg  _T_550; // @[package.scala 48:56:@39795.4]
  reg [31:0] _RAND_1;
  wire  x380_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x381_outr_UnitPipe.scala 101:55:@39801.4]
  wire  _T_563; // @[package.scala 96:25:@39828.4 package.scala 96:25:@39829.4]
  wire  _T_569; // @[package.scala 96:25:@39836.4 package.scala 96:25:@39837.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@39839.4]
  wire  x380_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@39840.4]
  x367_inr_UnitPipe_sm x367_inr_UnitPipe_sm ( // @[sm_x367_inr_UnitPipe.scala 33:18:@39319.4]
    .clock(x367_inr_UnitPipe_sm_clock),
    .reset(x367_inr_UnitPipe_sm_reset),
    .io_enable(x367_inr_UnitPipe_sm_io_enable),
    .io_done(x367_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x367_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x367_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x367_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x367_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x367_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x367_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39376.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39384.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1 x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1 ( // @[sm_x367_inr_UnitPipe.scala 69:24:@39414.4]
    .io_in_x360_valid(x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_valid),
    .io_in_x360_bits_addr(x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_bits_addr),
    .io_in_x360_bits_size(x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_bits_size),
    .io_in_x199_outdram_number(x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x199_outdram_number),
    .io_sigsIn_backpressure(x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_rr)
  );
  x369_ctrchain x369_ctrchain ( // @[SpatialBlocks.scala 37:22:@39482.4]
    .clock(x369_ctrchain_clock),
    .reset(x369_ctrchain_reset),
    .io_input_reset(x369_ctrchain_io_input_reset),
    .io_input_enable(x369_ctrchain_io_input_enable),
    .io_output_counts_0(x369_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x369_ctrchain_io_output_oobs_0),
    .io_output_done(x369_ctrchain_io_output_done)
  );
  x376_inr_Foreach_sm x376_inr_Foreach_sm ( // @[sm_x376_inr_Foreach.scala 33:18:@39535.4]
    .clock(x376_inr_Foreach_sm_clock),
    .reset(x376_inr_Foreach_sm_reset),
    .io_enable(x376_inr_Foreach_sm_io_enable),
    .io_done(x376_inr_Foreach_sm_io_done),
    .io_doneLatch(x376_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x376_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x376_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x376_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x376_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x376_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x376_inr_Foreach_sm_io_backpressure),
    .io_break(x376_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@39563.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@39603.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@39611.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x376_inr_Foreach_kernelx376_inr_Foreach_concrete1 x376_inr_Foreach_kernelx376_inr_Foreach_concrete1 ( // @[sm_x376_inr_Foreach.scala 78:24:@39646.4]
    .clock(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_clock),
    .reset(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_reset),
    .io_in_x361_valid(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_valid),
    .io_in_x361_bits_wdata_0(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_bits_wdata_0),
    .io_in_x361_bits_wstrb(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_bits_wstrb),
    .io_in_x203_outbuf_0_rPort_0_ofs_0(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0),
    .io_in_x203_outbuf_0_rPort_0_en_0(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_en_0),
    .io_in_x203_outbuf_0_rPort_0_backpressure(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure),
    .io_in_x203_outbuf_0_rPort_0_output_0(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_output_0),
    .io_sigsIn_backpressure(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_rr)
  );
  x380_inr_UnitPipe_sm x380_inr_UnitPipe_sm ( // @[sm_x380_inr_UnitPipe.scala 32:18:@39766.4]
    .clock(x380_inr_UnitPipe_sm_clock),
    .reset(x380_inr_UnitPipe_sm_reset),
    .io_enable(x380_inr_UnitPipe_sm_io_enable),
    .io_done(x380_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x380_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x380_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x380_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x380_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x380_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@39823.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@39831.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1 x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1 ( // @[sm_x380_inr_UnitPipe.scala 60:24:@39861.4]
    .io_in_x362_ready(x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1_io_in_x362_ready),
    .io_sigsIn_datapathEn(x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x367_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@39347.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@39381.4 package.scala 96:25:@39382.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@39389.4 package.scala 96:25:@39390.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@39392.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@39568.4 package.scala 96:25:@39569.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@39608.4 package.scala 96:25:@39609.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@39616.4 package.scala 96:25:@39617.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@39619.4]
  assign _T_479 = x376_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@39628.4]
  assign _T_480 = ~ x376_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@39629.4]
  assign _T_547 = x380_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@39794.4]
  assign x380_inr_UnitPipe_sigsIn_forwardpressure = io_in_x362_valid | x380_inr_UnitPipe_sm_io_doneLatch; // @[sm_x381_outr_UnitPipe.scala 101:55:@39801.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@39828.4 package.scala 96:25:@39829.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@39836.4 package.scala 96:25:@39837.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@39839.4]
  assign x380_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@39840.4]
  assign io_in_x361_valid = x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_valid; // @[sm_x376_inr_Foreach.scala 49:23:@39696.4]
  assign io_in_x361_bits_wdata_0 = x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_bits_wdata_0; // @[sm_x376_inr_Foreach.scala 49:23:@39695.4]
  assign io_in_x361_bits_wstrb = x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x361_bits_wstrb; // @[sm_x376_inr_Foreach.scala 49:23:@39694.4]
  assign io_in_x360_valid = x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_valid; // @[sm_x367_inr_UnitPipe.scala 49:23:@39452.4]
  assign io_in_x360_bits_addr = x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_bits_addr; // @[sm_x367_inr_UnitPipe.scala 49:23:@39451.4]
  assign io_in_x360_bits_size = x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x360_bits_size; // @[sm_x367_inr_UnitPipe.scala 49:23:@39450.4]
  assign io_in_x362_ready = x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1_io_in_x362_ready; // @[sm_x380_inr_UnitPipe.scala 46:23:@39897.4]
  assign io_in_x203_outbuf_0_rPort_0_ofs_0 = x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@39701.4]
  assign io_in_x203_outbuf_0_rPort_0_en_0 = x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@39700.4]
  assign io_in_x203_outbuf_0_rPort_0_backpressure = x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@39699.4]
  assign io_sigsOut_smDoneIn_0 = x367_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@39399.4]
  assign io_sigsOut_smDoneIn_1 = x376_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@39626.4]
  assign io_sigsOut_smDoneIn_2 = x380_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@39846.4]
  assign io_sigsOut_smCtrCopyDone_0 = x367_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@39413.4]
  assign io_sigsOut_smCtrCopyDone_1 = x376_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@39645.4]
  assign io_sigsOut_smCtrCopyDone_2 = x380_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@39860.4]
  assign x367_inr_UnitPipe_sm_clock = clock; // @[:@39320.4]
  assign x367_inr_UnitPipe_sm_reset = reset; // @[:@39321.4]
  assign x367_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@39396.4]
  assign x367_inr_UnitPipe_sm_io_ctrDone = x367_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x381_outr_UnitPipe.scala 77:39:@39351.4]
  assign x367_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@39398.4]
  assign x367_inr_UnitPipe_sm_io_backpressure = io_in_x360_ready | x367_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@39370.4]
  assign RetimeWrapper_clock = clock; // @[:@39377.4]
  assign RetimeWrapper_reset = reset; // @[:@39378.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39380.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@39379.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39385.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39386.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39388.4]
  assign RetimeWrapper_1_io_in = x367_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@39387.4]
  assign x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_in_x199_outdram_number = io_in_x199_outdram_number; // @[sm_x367_inr_UnitPipe.scala 50:31:@39454.4]
  assign x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x360_ready | x367_inr_UnitPipe_sm_io_doneLatch; // @[sm_x367_inr_UnitPipe.scala 74:22:@39469.4]
  assign x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x367_inr_UnitPipe_sm_io_datapathEn; // @[sm_x367_inr_UnitPipe.scala 74:22:@39467.4]
  assign x367_inr_UnitPipe_kernelx367_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x367_inr_UnitPipe.scala 73:18:@39455.4]
  assign x369_ctrchain_clock = clock; // @[:@39483.4]
  assign x369_ctrchain_reset = reset; // @[:@39484.4]
  assign x369_ctrchain_io_input_reset = x376_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@39644.4]
  assign x369_ctrchain_io_input_enable = x376_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@39596.4 SpatialBlocks.scala 159:42:@39643.4]
  assign x376_inr_Foreach_sm_clock = clock; // @[:@39536.4]
  assign x376_inr_Foreach_sm_reset = reset; // @[:@39537.4]
  assign x376_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@39623.4]
  assign x376_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x381_outr_UnitPipe.scala 90:38:@39571.4]
  assign x376_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@39625.4]
  assign x376_inr_Foreach_sm_io_backpressure = io_in_x361_ready | x376_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@39597.4]
  assign x376_inr_Foreach_sm_io_break = 1'h0; // @[sm_x381_outr_UnitPipe.scala 94:36:@39577.4]
  assign RetimeWrapper_2_clock = clock; // @[:@39564.4]
  assign RetimeWrapper_2_reset = reset; // @[:@39565.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@39567.4]
  assign RetimeWrapper_2_io_in = x369_ctrchain_io_output_done; // @[package.scala 94:16:@39566.4]
  assign RetimeWrapper_3_clock = clock; // @[:@39604.4]
  assign RetimeWrapper_3_reset = reset; // @[:@39605.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@39607.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@39606.4]
  assign RetimeWrapper_4_clock = clock; // @[:@39612.4]
  assign RetimeWrapper_4_reset = reset; // @[:@39613.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@39615.4]
  assign RetimeWrapper_4_io_in = x376_inr_Foreach_sm_io_done; // @[package.scala 94:16:@39614.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_clock = clock; // @[:@39647.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_reset = reset; // @[:@39648.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_in_x203_outbuf_0_rPort_0_output_0 = io_in_x203_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@39698.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x361_ready | x376_inr_Foreach_sm_io_doneLatch; // @[sm_x376_inr_Foreach.scala 83:22:@39717.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x376_inr_Foreach.scala 83:22:@39715.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_break = x376_inr_Foreach_sm_io_break; // @[sm_x376_inr_Foreach.scala 83:22:@39713.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x369_ctrchain_io_output_counts_0[22]}},x369_ctrchain_io_output_counts_0}; // @[sm_x376_inr_Foreach.scala 83:22:@39708.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x369_ctrchain_io_output_oobs_0; // @[sm_x376_inr_Foreach.scala 83:22:@39707.4]
  assign x376_inr_Foreach_kernelx376_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x376_inr_Foreach.scala 82:18:@39703.4]
  assign x380_inr_UnitPipe_sm_clock = clock; // @[:@39767.4]
  assign x380_inr_UnitPipe_sm_reset = reset; // @[:@39768.4]
  assign x380_inr_UnitPipe_sm_io_enable = x380_inr_UnitPipe_sigsIn_baseEn & x380_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@39843.4]
  assign x380_inr_UnitPipe_sm_io_ctrDone = x380_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x381_outr_UnitPipe.scala 99:39:@39798.4]
  assign x380_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@39845.4]
  assign RetimeWrapper_5_clock = clock; // @[:@39824.4]
  assign RetimeWrapper_5_reset = reset; // @[:@39825.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@39827.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@39826.4]
  assign RetimeWrapper_6_clock = clock; // @[:@39832.4]
  assign RetimeWrapper_6_reset = reset; // @[:@39833.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@39835.4]
  assign RetimeWrapper_6_io_in = x380_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@39834.4]
  assign x380_inr_UnitPipe_kernelx380_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x380_inr_UnitPipe_sm_io_datapathEn; // @[sm_x380_inr_UnitPipe.scala 65:22:@39910.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x491_kernelx491_concrete1( // @[:@39926.2]
  input          clock, // @[:@39927.4]
  input          reset, // @[:@39928.4]
  output         io_in_x202_TVALID, // @[:@39929.4]
  input          io_in_x202_TREADY, // @[:@39929.4]
  output [255:0] io_in_x202_TDATA, // @[:@39929.4]
  input          io_in_x201_TVALID, // @[:@39929.4]
  output         io_in_x201_TREADY, // @[:@39929.4]
  input  [255:0] io_in_x201_TDATA, // @[:@39929.4]
  input  [7:0]   io_in_x201_TID, // @[:@39929.4]
  input  [7:0]   io_in_x201_TDEST, // @[:@39929.4]
  input          io_in_x361_ready, // @[:@39929.4]
  output         io_in_x361_valid, // @[:@39929.4]
  output [31:0]  io_in_x361_bits_wdata_0, // @[:@39929.4]
  output         io_in_x361_bits_wstrb, // @[:@39929.4]
  input          io_in_x360_ready, // @[:@39929.4]
  output         io_in_x360_valid, // @[:@39929.4]
  output [63:0]  io_in_x360_bits_addr, // @[:@39929.4]
  output [31:0]  io_in_x360_bits_size, // @[:@39929.4]
  output         io_in_x362_ready, // @[:@39929.4]
  input          io_in_x362_valid, // @[:@39929.4]
  input  [63:0]  io_in_x199_outdram_number, // @[:@39929.4]
  output [20:0]  io_in_x203_outbuf_0_rPort_0_ofs_0, // @[:@39929.4]
  output         io_in_x203_outbuf_0_rPort_0_en_0, // @[:@39929.4]
  output         io_in_x203_outbuf_0_rPort_0_backpressure, // @[:@39929.4]
  input  [31:0]  io_in_x203_outbuf_0_rPort_0_output_0, // @[:@39929.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@39929.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@39929.4]
  input          io_sigsIn_smChildAcks_0, // @[:@39929.4]
  input          io_sigsIn_smChildAcks_1, // @[:@39929.4]
  output         io_sigsOut_smDoneIn_0, // @[:@39929.4]
  output         io_sigsOut_smDoneIn_1, // @[:@39929.4]
  input          io_rr // @[:@39929.4]
);
  wire  x359_outr_UnitPipe_sm_clock; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_reset; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_enable; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_done; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_parentAck; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_childAck_0; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_childAck_1; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  x359_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@40064.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@40064.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@40064.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@40064.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@40064.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@40072.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@40072.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@40072.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@40072.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@40072.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_clock; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_reset; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TVALID; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TREADY; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire [255:0] x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TDATA; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TVALID; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TREADY; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire [255:0] x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TDATA; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire [7:0] x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TID; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire [7:0] x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TDEST; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_rr; // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
  wire  x381_outr_UnitPipe_sm_clock; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_reset; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_enable; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_done; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_parentAck; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_childAck_0; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_childAck_1; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_childAck_2; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  x381_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@40353.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@40353.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@40353.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@40353.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@40353.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@40361.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@40361.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@40361.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@40361.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@40361.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_clock; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_reset; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_ready; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_valid; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire [31:0] x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_bits_wdata_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_bits_wstrb; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_ready; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_valid; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire [63:0] x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_bits_addr; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire [31:0] x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_bits_size; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x362_ready; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x362_valid; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire [63:0] x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x199_outdram_number; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire [20:0] x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_en_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire [31:0] x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_output_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_rr; // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
  wire  _T_408; // @[package.scala 96:25:@40069.4 package.scala 96:25:@40070.4]
  wire  _T_414; // @[package.scala 96:25:@40077.4 package.scala 96:25:@40078.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@40080.4]
  wire  _T_508; // @[package.scala 96:25:@40358.4 package.scala 96:25:@40359.4]
  wire  _T_514; // @[package.scala 96:25:@40366.4 package.scala 96:25:@40367.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@40369.4]
  x359_outr_UnitPipe_sm x359_outr_UnitPipe_sm ( // @[sm_x359_outr_UnitPipe.scala 32:18:@40002.4]
    .clock(x359_outr_UnitPipe_sm_clock),
    .reset(x359_outr_UnitPipe_sm_reset),
    .io_enable(x359_outr_UnitPipe_sm_io_enable),
    .io_done(x359_outr_UnitPipe_sm_io_done),
    .io_parentAck(x359_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x359_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x359_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x359_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x359_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x359_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x359_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x359_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x359_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@40064.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@40072.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1 x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1 ( // @[sm_x359_outr_UnitPipe.scala 87:24:@40103.4]
    .clock(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_clock),
    .reset(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_reset),
    .io_in_x202_TVALID(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TVALID),
    .io_in_x202_TREADY(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TREADY),
    .io_in_x202_TDATA(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TDATA),
    .io_in_x201_TVALID(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TVALID),
    .io_in_x201_TREADY(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TREADY),
    .io_in_x201_TDATA(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TDATA),
    .io_in_x201_TID(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TID),
    .io_in_x201_TDEST(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TDEST),
    .io_sigsIn_smEnableOuts_0(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_rr)
  );
  x381_outr_UnitPipe_sm x381_outr_UnitPipe_sm ( // @[sm_x381_outr_UnitPipe.scala 36:18:@40281.4]
    .clock(x381_outr_UnitPipe_sm_clock),
    .reset(x381_outr_UnitPipe_sm_reset),
    .io_enable(x381_outr_UnitPipe_sm_io_enable),
    .io_done(x381_outr_UnitPipe_sm_io_done),
    .io_parentAck(x381_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x381_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x381_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x381_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x381_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x381_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x381_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x381_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x381_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x381_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x381_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x381_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x381_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@40353.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@40361.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1 x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1 ( // @[sm_x381_outr_UnitPipe.scala 108:24:@40393.4]
    .clock(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_clock),
    .reset(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_reset),
    .io_in_x361_ready(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_ready),
    .io_in_x361_valid(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_valid),
    .io_in_x361_bits_wdata_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_bits_wdata_0),
    .io_in_x361_bits_wstrb(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_bits_wstrb),
    .io_in_x360_ready(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_ready),
    .io_in_x360_valid(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_valid),
    .io_in_x360_bits_addr(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_bits_addr),
    .io_in_x360_bits_size(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_bits_size),
    .io_in_x362_ready(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x362_ready),
    .io_in_x362_valid(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x362_valid),
    .io_in_x199_outdram_number(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x199_outdram_number),
    .io_in_x203_outbuf_0_rPort_0_ofs_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0),
    .io_in_x203_outbuf_0_rPort_0_en_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_en_0),
    .io_in_x203_outbuf_0_rPort_0_backpressure(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure),
    .io_in_x203_outbuf_0_rPort_0_output_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_output_0),
    .io_sigsIn_smEnableOuts_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@40069.4 package.scala 96:25:@40070.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@40077.4 package.scala 96:25:@40078.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@40080.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@40358.4 package.scala 96:25:@40359.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@40366.4 package.scala 96:25:@40367.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@40369.4]
  assign io_in_x202_TVALID = x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TVALID; // @[sm_x359_outr_UnitPipe.scala 48:23:@40172.4]
  assign io_in_x202_TDATA = x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TDATA; // @[sm_x359_outr_UnitPipe.scala 48:23:@40170.4]
  assign io_in_x201_TREADY = x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TREADY; // @[sm_x359_outr_UnitPipe.scala 49:23:@40180.4]
  assign io_in_x361_valid = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_valid; // @[sm_x381_outr_UnitPipe.scala 58:23:@40475.4]
  assign io_in_x361_bits_wdata_0 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_bits_wdata_0; // @[sm_x381_outr_UnitPipe.scala 58:23:@40474.4]
  assign io_in_x361_bits_wstrb = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_bits_wstrb; // @[sm_x381_outr_UnitPipe.scala 58:23:@40473.4]
  assign io_in_x360_valid = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_valid; // @[sm_x381_outr_UnitPipe.scala 59:23:@40479.4]
  assign io_in_x360_bits_addr = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_bits_addr; // @[sm_x381_outr_UnitPipe.scala 59:23:@40478.4]
  assign io_in_x360_bits_size = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_bits_size; // @[sm_x381_outr_UnitPipe.scala 59:23:@40477.4]
  assign io_in_x362_ready = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x362_ready; // @[sm_x381_outr_UnitPipe.scala 60:23:@40483.4]
  assign io_in_x203_outbuf_0_rPort_0_ofs_0 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@40488.4]
  assign io_in_x203_outbuf_0_rPort_0_en_0 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@40487.4]
  assign io_in_x203_outbuf_0_rPort_0_backpressure = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@40486.4]
  assign io_sigsOut_smDoneIn_0 = x359_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@40087.4]
  assign io_sigsOut_smDoneIn_1 = x381_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@40376.4]
  assign x359_outr_UnitPipe_sm_clock = clock; // @[:@40003.4]
  assign x359_outr_UnitPipe_sm_reset = reset; // @[:@40004.4]
  assign x359_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@40084.4]
  assign x359_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@40086.4]
  assign x359_outr_UnitPipe_sm_io_doneIn_0 = x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@40054.4]
  assign x359_outr_UnitPipe_sm_io_doneIn_1 = x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@40055.4]
  assign x359_outr_UnitPipe_sm_io_ctrCopyDone_0 = x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@40101.4]
  assign x359_outr_UnitPipe_sm_io_ctrCopyDone_1 = x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@40102.4]
  assign RetimeWrapper_clock = clock; // @[:@40065.4]
  assign RetimeWrapper_reset = reset; // @[:@40066.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@40068.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@40067.4]
  assign RetimeWrapper_1_clock = clock; // @[:@40073.4]
  assign RetimeWrapper_1_reset = reset; // @[:@40074.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@40076.4]
  assign RetimeWrapper_1_io_in = x359_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@40075.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_clock = clock; // @[:@40104.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_reset = reset; // @[:@40105.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x202_TREADY = io_in_x202_TREADY; // @[sm_x359_outr_UnitPipe.scala 48:23:@40171.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TVALID = io_in_x201_TVALID; // @[sm_x359_outr_UnitPipe.scala 49:23:@40181.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TDATA = io_in_x201_TDATA; // @[sm_x359_outr_UnitPipe.scala 49:23:@40179.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TID = io_in_x201_TID; // @[sm_x359_outr_UnitPipe.scala 49:23:@40175.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_in_x201_TDEST = io_in_x201_TDEST; // @[sm_x359_outr_UnitPipe.scala 49:23:@40174.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x359_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x359_outr_UnitPipe.scala 92:22:@40197.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x359_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x359_outr_UnitPipe.scala 92:22:@40198.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x359_outr_UnitPipe_sm_io_childAck_0; // @[sm_x359_outr_UnitPipe.scala 92:22:@40193.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x359_outr_UnitPipe_sm_io_childAck_1; // @[sm_x359_outr_UnitPipe.scala 92:22:@40194.4]
  assign x359_outr_UnitPipe_kernelx359_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x359_outr_UnitPipe.scala 91:18:@40182.4]
  assign x381_outr_UnitPipe_sm_clock = clock; // @[:@40282.4]
  assign x381_outr_UnitPipe_sm_reset = reset; // @[:@40283.4]
  assign x381_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@40373.4]
  assign x381_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@40375.4]
  assign x381_outr_UnitPipe_sm_io_doneIn_0 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@40341.4]
  assign x381_outr_UnitPipe_sm_io_doneIn_1 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@40342.4]
  assign x381_outr_UnitPipe_sm_io_doneIn_2 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@40343.4]
  assign x381_outr_UnitPipe_sm_io_ctrCopyDone_0 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@40390.4]
  assign x381_outr_UnitPipe_sm_io_ctrCopyDone_1 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@40391.4]
  assign x381_outr_UnitPipe_sm_io_ctrCopyDone_2 = x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@40392.4]
  assign RetimeWrapper_2_clock = clock; // @[:@40354.4]
  assign RetimeWrapper_2_reset = reset; // @[:@40355.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@40357.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@40356.4]
  assign RetimeWrapper_3_clock = clock; // @[:@40362.4]
  assign RetimeWrapper_3_reset = reset; // @[:@40363.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@40365.4]
  assign RetimeWrapper_3_io_in = x381_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@40364.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_clock = clock; // @[:@40394.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_reset = reset; // @[:@40395.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x361_ready = io_in_x361_ready; // @[sm_x381_outr_UnitPipe.scala 58:23:@40476.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x360_ready = io_in_x360_ready; // @[sm_x381_outr_UnitPipe.scala 59:23:@40480.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x362_valid = io_in_x362_valid; // @[sm_x381_outr_UnitPipe.scala 60:23:@40482.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x199_outdram_number = io_in_x199_outdram_number; // @[sm_x381_outr_UnitPipe.scala 61:31:@40484.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_in_x203_outbuf_0_rPort_0_output_0 = io_in_x203_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@40485.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x381_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x381_outr_UnitPipe.scala 113:22:@40512.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x381_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x381_outr_UnitPipe.scala 113:22:@40513.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x381_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x381_outr_UnitPipe.scala 113:22:@40514.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x381_outr_UnitPipe_sm_io_childAck_0; // @[sm_x381_outr_UnitPipe.scala 113:22:@40506.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x381_outr_UnitPipe_sm_io_childAck_1; // @[sm_x381_outr_UnitPipe.scala 113:22:@40507.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x381_outr_UnitPipe_sm_io_childAck_2; // @[sm_x381_outr_UnitPipe.scala 113:22:@40508.4]
  assign x381_outr_UnitPipe_kernelx381_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x381_outr_UnitPipe.scala 112:18:@40490.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@40542.2]
  input          clock, // @[:@40543.4]
  input          reset, // @[:@40544.4]
  output         io_in_x202_TVALID, // @[:@40545.4]
  input          io_in_x202_TREADY, // @[:@40545.4]
  output [255:0] io_in_x202_TDATA, // @[:@40545.4]
  input          io_in_x201_TVALID, // @[:@40545.4]
  output         io_in_x201_TREADY, // @[:@40545.4]
  input  [255:0] io_in_x201_TDATA, // @[:@40545.4]
  input  [7:0]   io_in_x201_TID, // @[:@40545.4]
  input  [7:0]   io_in_x201_TDEST, // @[:@40545.4]
  input          io_in_x361_ready, // @[:@40545.4]
  output         io_in_x361_valid, // @[:@40545.4]
  output [31:0]  io_in_x361_bits_wdata_0, // @[:@40545.4]
  output         io_in_x361_bits_wstrb, // @[:@40545.4]
  input          io_in_x360_ready, // @[:@40545.4]
  output         io_in_x360_valid, // @[:@40545.4]
  output [63:0]  io_in_x360_bits_addr, // @[:@40545.4]
  output [31:0]  io_in_x360_bits_size, // @[:@40545.4]
  output         io_in_x362_ready, // @[:@40545.4]
  input          io_in_x362_valid, // @[:@40545.4]
  input  [63:0]  io_in_x199_outdram_number, // @[:@40545.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@40545.4]
  input          io_sigsIn_smChildAcks_0, // @[:@40545.4]
  output         io_sigsOut_smDoneIn_0, // @[:@40545.4]
  input          io_rr // @[:@40545.4]
);
  wire  x203_outbuf_0_clock; // @[m_x203_outbuf_0.scala 27:17:@40555.4]
  wire  x203_outbuf_0_reset; // @[m_x203_outbuf_0.scala 27:17:@40555.4]
  wire [20:0] x203_outbuf_0_io_rPort_0_ofs_0; // @[m_x203_outbuf_0.scala 27:17:@40555.4]
  wire  x203_outbuf_0_io_rPort_0_en_0; // @[m_x203_outbuf_0.scala 27:17:@40555.4]
  wire  x203_outbuf_0_io_rPort_0_backpressure; // @[m_x203_outbuf_0.scala 27:17:@40555.4]
  wire [31:0] x203_outbuf_0_io_rPort_0_output_0; // @[m_x203_outbuf_0.scala 27:17:@40555.4]
  wire  x491_sm_clock; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_reset; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_enable; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_done; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_ctrDone; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_ctrInc; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_parentAck; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_doneIn_0; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_doneIn_1; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_enableOut_0; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_enableOut_1; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_childAck_0; // @[sm_x491.scala 37:18:@40613.4]
  wire  x491_sm_io_childAck_1; // @[sm_x491.scala 37:18:@40613.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@40680.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@40680.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@40680.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@40680.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@40680.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@40688.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@40688.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@40688.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@40688.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@40688.4]
  wire  x491_kernelx491_concrete1_clock; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_reset; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x202_TVALID; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x202_TREADY; // @[sm_x491.scala 102:24:@40717.4]
  wire [255:0] x491_kernelx491_concrete1_io_in_x202_TDATA; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x201_TVALID; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x201_TREADY; // @[sm_x491.scala 102:24:@40717.4]
  wire [255:0] x491_kernelx491_concrete1_io_in_x201_TDATA; // @[sm_x491.scala 102:24:@40717.4]
  wire [7:0] x491_kernelx491_concrete1_io_in_x201_TID; // @[sm_x491.scala 102:24:@40717.4]
  wire [7:0] x491_kernelx491_concrete1_io_in_x201_TDEST; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x361_ready; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x361_valid; // @[sm_x491.scala 102:24:@40717.4]
  wire [31:0] x491_kernelx491_concrete1_io_in_x361_bits_wdata_0; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x361_bits_wstrb; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x360_ready; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x360_valid; // @[sm_x491.scala 102:24:@40717.4]
  wire [63:0] x491_kernelx491_concrete1_io_in_x360_bits_addr; // @[sm_x491.scala 102:24:@40717.4]
  wire [31:0] x491_kernelx491_concrete1_io_in_x360_bits_size; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x362_ready; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x362_valid; // @[sm_x491.scala 102:24:@40717.4]
  wire [63:0] x491_kernelx491_concrete1_io_in_x199_outdram_number; // @[sm_x491.scala 102:24:@40717.4]
  wire [20:0] x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_en_0; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure; // @[sm_x491.scala 102:24:@40717.4]
  wire [31:0] x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_output_0; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x491.scala 102:24:@40717.4]
  wire  x491_kernelx491_concrete1_io_rr; // @[sm_x491.scala 102:24:@40717.4]
  wire  _T_266; // @[package.scala 100:49:@40646.4]
  reg  _T_269; // @[package.scala 48:56:@40647.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@40685.4 package.scala 96:25:@40686.4]
  wire  _T_289; // @[package.scala 96:25:@40693.4 package.scala 96:25:@40694.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@40696.4]
  x203_outbuf_0 x203_outbuf_0 ( // @[m_x203_outbuf_0.scala 27:17:@40555.4]
    .clock(x203_outbuf_0_clock),
    .reset(x203_outbuf_0_reset),
    .io_rPort_0_ofs_0(x203_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x203_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x203_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x203_outbuf_0_io_rPort_0_output_0)
  );
  x491_sm x491_sm ( // @[sm_x491.scala 37:18:@40613.4]
    .clock(x491_sm_clock),
    .reset(x491_sm_reset),
    .io_enable(x491_sm_io_enable),
    .io_done(x491_sm_io_done),
    .io_ctrDone(x491_sm_io_ctrDone),
    .io_ctrInc(x491_sm_io_ctrInc),
    .io_parentAck(x491_sm_io_parentAck),
    .io_doneIn_0(x491_sm_io_doneIn_0),
    .io_doneIn_1(x491_sm_io_doneIn_1),
    .io_enableOut_0(x491_sm_io_enableOut_0),
    .io_enableOut_1(x491_sm_io_enableOut_1),
    .io_childAck_0(x491_sm_io_childAck_0),
    .io_childAck_1(x491_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@40680.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@40688.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x491_kernelx491_concrete1 x491_kernelx491_concrete1 ( // @[sm_x491.scala 102:24:@40717.4]
    .clock(x491_kernelx491_concrete1_clock),
    .reset(x491_kernelx491_concrete1_reset),
    .io_in_x202_TVALID(x491_kernelx491_concrete1_io_in_x202_TVALID),
    .io_in_x202_TREADY(x491_kernelx491_concrete1_io_in_x202_TREADY),
    .io_in_x202_TDATA(x491_kernelx491_concrete1_io_in_x202_TDATA),
    .io_in_x201_TVALID(x491_kernelx491_concrete1_io_in_x201_TVALID),
    .io_in_x201_TREADY(x491_kernelx491_concrete1_io_in_x201_TREADY),
    .io_in_x201_TDATA(x491_kernelx491_concrete1_io_in_x201_TDATA),
    .io_in_x201_TID(x491_kernelx491_concrete1_io_in_x201_TID),
    .io_in_x201_TDEST(x491_kernelx491_concrete1_io_in_x201_TDEST),
    .io_in_x361_ready(x491_kernelx491_concrete1_io_in_x361_ready),
    .io_in_x361_valid(x491_kernelx491_concrete1_io_in_x361_valid),
    .io_in_x361_bits_wdata_0(x491_kernelx491_concrete1_io_in_x361_bits_wdata_0),
    .io_in_x361_bits_wstrb(x491_kernelx491_concrete1_io_in_x361_bits_wstrb),
    .io_in_x360_ready(x491_kernelx491_concrete1_io_in_x360_ready),
    .io_in_x360_valid(x491_kernelx491_concrete1_io_in_x360_valid),
    .io_in_x360_bits_addr(x491_kernelx491_concrete1_io_in_x360_bits_addr),
    .io_in_x360_bits_size(x491_kernelx491_concrete1_io_in_x360_bits_size),
    .io_in_x362_ready(x491_kernelx491_concrete1_io_in_x362_ready),
    .io_in_x362_valid(x491_kernelx491_concrete1_io_in_x362_valid),
    .io_in_x199_outdram_number(x491_kernelx491_concrete1_io_in_x199_outdram_number),
    .io_in_x203_outbuf_0_rPort_0_ofs_0(x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0),
    .io_in_x203_outbuf_0_rPort_0_en_0(x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_en_0),
    .io_in_x203_outbuf_0_rPort_0_backpressure(x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure),
    .io_in_x203_outbuf_0_rPort_0_output_0(x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_output_0),
    .io_sigsIn_smEnableOuts_0(x491_kernelx491_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x491_kernelx491_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x491_kernelx491_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x491_kernelx491_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x491_kernelx491_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x491_kernelx491_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x491_kernelx491_concrete1_io_rr)
  );
  assign _T_266 = x491_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@40646.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@40685.4 package.scala 96:25:@40686.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@40693.4 package.scala 96:25:@40694.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@40696.4]
  assign io_in_x202_TVALID = x491_kernelx491_concrete1_io_in_x202_TVALID; // @[sm_x491.scala 63:23:@40804.4]
  assign io_in_x202_TDATA = x491_kernelx491_concrete1_io_in_x202_TDATA; // @[sm_x491.scala 63:23:@40802.4]
  assign io_in_x201_TREADY = x491_kernelx491_concrete1_io_in_x201_TREADY; // @[sm_x491.scala 64:23:@40812.4]
  assign io_in_x361_valid = x491_kernelx491_concrete1_io_in_x361_valid; // @[sm_x491.scala 65:23:@40816.4]
  assign io_in_x361_bits_wdata_0 = x491_kernelx491_concrete1_io_in_x361_bits_wdata_0; // @[sm_x491.scala 65:23:@40815.4]
  assign io_in_x361_bits_wstrb = x491_kernelx491_concrete1_io_in_x361_bits_wstrb; // @[sm_x491.scala 65:23:@40814.4]
  assign io_in_x360_valid = x491_kernelx491_concrete1_io_in_x360_valid; // @[sm_x491.scala 66:23:@40820.4]
  assign io_in_x360_bits_addr = x491_kernelx491_concrete1_io_in_x360_bits_addr; // @[sm_x491.scala 66:23:@40819.4]
  assign io_in_x360_bits_size = x491_kernelx491_concrete1_io_in_x360_bits_size; // @[sm_x491.scala 66:23:@40818.4]
  assign io_in_x362_ready = x491_kernelx491_concrete1_io_in_x362_ready; // @[sm_x491.scala 67:23:@40824.4]
  assign io_sigsOut_smDoneIn_0 = x491_sm_io_done; // @[SpatialBlocks.scala 156:53:@40703.4]
  assign x203_outbuf_0_clock = clock; // @[:@40556.4]
  assign x203_outbuf_0_reset = reset; // @[:@40557.4]
  assign x203_outbuf_0_io_rPort_0_ofs_0 = x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@40829.4]
  assign x203_outbuf_0_io_rPort_0_en_0 = x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@40828.4]
  assign x203_outbuf_0_io_rPort_0_backpressure = x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@40827.4]
  assign x491_sm_clock = clock; // @[:@40614.4]
  assign x491_sm_reset = reset; // @[:@40615.4]
  assign x491_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@40700.4]
  assign x491_sm_io_ctrDone = x491_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@40650.4]
  assign x491_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@40702.4]
  assign x491_sm_io_doneIn_0 = x491_kernelx491_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@40670.4]
  assign x491_sm_io_doneIn_1 = x491_kernelx491_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@40671.4]
  assign RetimeWrapper_clock = clock; // @[:@40681.4]
  assign RetimeWrapper_reset = reset; // @[:@40682.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@40684.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@40683.4]
  assign RetimeWrapper_1_clock = clock; // @[:@40689.4]
  assign RetimeWrapper_1_reset = reset; // @[:@40690.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@40692.4]
  assign RetimeWrapper_1_io_in = x491_sm_io_done; // @[package.scala 94:16:@40691.4]
  assign x491_kernelx491_concrete1_clock = clock; // @[:@40718.4]
  assign x491_kernelx491_concrete1_reset = reset; // @[:@40719.4]
  assign x491_kernelx491_concrete1_io_in_x202_TREADY = io_in_x202_TREADY; // @[sm_x491.scala 63:23:@40803.4]
  assign x491_kernelx491_concrete1_io_in_x201_TVALID = io_in_x201_TVALID; // @[sm_x491.scala 64:23:@40813.4]
  assign x491_kernelx491_concrete1_io_in_x201_TDATA = io_in_x201_TDATA; // @[sm_x491.scala 64:23:@40811.4]
  assign x491_kernelx491_concrete1_io_in_x201_TID = io_in_x201_TID; // @[sm_x491.scala 64:23:@40807.4]
  assign x491_kernelx491_concrete1_io_in_x201_TDEST = io_in_x201_TDEST; // @[sm_x491.scala 64:23:@40806.4]
  assign x491_kernelx491_concrete1_io_in_x361_ready = io_in_x361_ready; // @[sm_x491.scala 65:23:@40817.4]
  assign x491_kernelx491_concrete1_io_in_x360_ready = io_in_x360_ready; // @[sm_x491.scala 66:23:@40821.4]
  assign x491_kernelx491_concrete1_io_in_x362_valid = io_in_x362_valid; // @[sm_x491.scala 67:23:@40823.4]
  assign x491_kernelx491_concrete1_io_in_x199_outdram_number = io_in_x199_outdram_number; // @[sm_x491.scala 68:31:@40825.4]
  assign x491_kernelx491_concrete1_io_in_x203_outbuf_0_rPort_0_output_0 = x203_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@40826.4]
  assign x491_kernelx491_concrete1_io_sigsIn_smEnableOuts_0 = x491_sm_io_enableOut_0; // @[sm_x491.scala 107:22:@40841.4]
  assign x491_kernelx491_concrete1_io_sigsIn_smEnableOuts_1 = x491_sm_io_enableOut_1; // @[sm_x491.scala 107:22:@40842.4]
  assign x491_kernelx491_concrete1_io_sigsIn_smChildAcks_0 = x491_sm_io_childAck_0; // @[sm_x491.scala 107:22:@40837.4]
  assign x491_kernelx491_concrete1_io_sigsIn_smChildAcks_1 = x491_sm_io_childAck_1; // @[sm_x491.scala 107:22:@40838.4]
  assign x491_kernelx491_concrete1_io_rr = io_rr; // @[sm_x491.scala 106:18:@40831.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@40864.2]
  input          clock, // @[:@40865.4]
  input          reset, // @[:@40866.4]
  input          io_enable, // @[:@40867.4]
  output         io_done, // @[:@40867.4]
  input          io_reset, // @[:@40867.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@40867.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@40867.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@40867.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@40867.4]
  output         io_memStreams_loads_0_data_ready, // @[:@40867.4]
  input          io_memStreams_loads_0_data_valid, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@40867.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@40867.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@40867.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@40867.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@40867.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@40867.4]
  input          io_memStreams_stores_0_data_ready, // @[:@40867.4]
  output         io_memStreams_stores_0_data_valid, // @[:@40867.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@40867.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@40867.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@40867.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@40867.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@40867.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@40867.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@40867.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@40867.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@40867.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@40867.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@40867.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@40867.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@40867.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@40867.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@40867.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@40867.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@40867.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@40867.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@40867.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@40867.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@40867.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@40867.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@40867.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@40867.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@40867.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@40867.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@40867.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@40867.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@40867.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@40867.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@40867.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@40867.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@40867.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@40867.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@40867.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@40867.4]
  output         io_heap_0_req_valid, // @[:@40867.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@40867.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@40867.4]
  input          io_heap_0_resp_valid, // @[:@40867.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@40867.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@40867.4]
  input  [63:0]  io_argIns_0, // @[:@40867.4]
  input  [63:0]  io_argIns_1, // @[:@40867.4]
  input          io_argOuts_0_port_ready, // @[:@40867.4]
  output         io_argOuts_0_port_valid, // @[:@40867.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@40867.4]
  input  [63:0]  io_argOuts_0_echo // @[:@40867.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@41015.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@41015.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@41015.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@41015.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41033.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41033.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41033.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@41033.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@41033.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@41042.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@41042.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@41042.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@41042.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@41042.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@41042.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@41081.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@41113.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@41113.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@41113.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@41113.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@41113.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x202_TVALID; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x202_TREADY; // @[sm_RootController.scala 91:24:@41175.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x202_TDATA; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x201_TVALID; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x201_TREADY; // @[sm_RootController.scala 91:24:@41175.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x201_TDATA; // @[sm_RootController.scala 91:24:@41175.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x201_TID; // @[sm_RootController.scala 91:24:@41175.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x201_TDEST; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x361_ready; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x361_valid; // @[sm_RootController.scala 91:24:@41175.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x361_bits_wdata_0; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x361_bits_wstrb; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x360_ready; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x360_valid; // @[sm_RootController.scala 91:24:@41175.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x360_bits_addr; // @[sm_RootController.scala 91:24:@41175.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x360_bits_size; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x362_ready; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_in_x362_valid; // @[sm_RootController.scala 91:24:@41175.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x199_outdram_number; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@41175.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@41175.4]
  wire  _T_599; // @[package.scala 96:25:@41038.4 package.scala 96:25:@41039.4]
  wire  _T_664; // @[Main.scala 46:50:@41109.4]
  wire  _T_665; // @[Main.scala 46:59:@41110.4]
  wire  _T_677; // @[package.scala 100:49:@41130.4]
  reg  _T_680; // @[package.scala 48:56:@41131.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@41015.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@41033.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@41042.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@41081.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@41113.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@41175.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x202_TVALID(RootController_kernelRootController_concrete1_io_in_x202_TVALID),
    .io_in_x202_TREADY(RootController_kernelRootController_concrete1_io_in_x202_TREADY),
    .io_in_x202_TDATA(RootController_kernelRootController_concrete1_io_in_x202_TDATA),
    .io_in_x201_TVALID(RootController_kernelRootController_concrete1_io_in_x201_TVALID),
    .io_in_x201_TREADY(RootController_kernelRootController_concrete1_io_in_x201_TREADY),
    .io_in_x201_TDATA(RootController_kernelRootController_concrete1_io_in_x201_TDATA),
    .io_in_x201_TID(RootController_kernelRootController_concrete1_io_in_x201_TID),
    .io_in_x201_TDEST(RootController_kernelRootController_concrete1_io_in_x201_TDEST),
    .io_in_x361_ready(RootController_kernelRootController_concrete1_io_in_x361_ready),
    .io_in_x361_valid(RootController_kernelRootController_concrete1_io_in_x361_valid),
    .io_in_x361_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x361_bits_wdata_0),
    .io_in_x361_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x361_bits_wstrb),
    .io_in_x360_ready(RootController_kernelRootController_concrete1_io_in_x360_ready),
    .io_in_x360_valid(RootController_kernelRootController_concrete1_io_in_x360_valid),
    .io_in_x360_bits_addr(RootController_kernelRootController_concrete1_io_in_x360_bits_addr),
    .io_in_x360_bits_size(RootController_kernelRootController_concrete1_io_in_x360_bits_size),
    .io_in_x362_ready(RootController_kernelRootController_concrete1_io_in_x362_ready),
    .io_in_x362_valid(RootController_kernelRootController_concrete1_io_in_x362_valid),
    .io_in_x199_outdram_number(RootController_kernelRootController_concrete1_io_in_x199_outdram_number),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@41038.4 package.scala 96:25:@41039.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@41109.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@41110.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@41130.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@41129.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x360_valid; // @[sm_RootController.scala 63:23:@41260.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x360_bits_addr; // @[sm_RootController.scala 63:23:@41259.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x360_bits_size; // @[sm_RootController.scala 63:23:@41258.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x361_valid; // @[sm_RootController.scala 62:23:@41256.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x361_bits_wdata_0; // @[sm_RootController.scala 62:23:@41255.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x361_bits_wstrb; // @[sm_RootController.scala 62:23:@41254.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x362_ready; // @[sm_RootController.scala 64:23:@41264.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x201_TREADY; // @[sm_RootController.scala 61:23:@41252.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x202_TVALID; // @[sm_RootController.scala 60:23:@41244.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x202_TDATA; // @[sm_RootController.scala 60:23:@41242.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 60:23:@41241.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 60:23:@41240.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 60:23:@41239.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 60:23:@41238.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 60:23:@41237.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 60:23:@41236.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@41016.4]
  assign SingleCounter_reset = reset; // @[:@41017.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@41031.4]
  assign RetimeWrapper_clock = clock; // @[:@41034.4]
  assign RetimeWrapper_reset = reset; // @[:@41035.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@41037.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@41036.4]
  assign SRFF_clock = clock; // @[:@41043.4]
  assign SRFF_reset = reset; // @[:@41044.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@41293.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@41127.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@41128.4]
  assign RootController_sm_clock = clock; // @[:@41082.4]
  assign RootController_sm_reset = reset; // @[:@41083.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@41126.4 SpatialBlocks.scala 140:18:@41160.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@41154.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@41134.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@41122.4 SpatialBlocks.scala 142:21:@41162.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@41151.4]
  assign RetimeWrapper_1_clock = clock; // @[:@41114.4]
  assign RetimeWrapper_1_reset = reset; // @[:@41115.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@41117.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@41116.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@41176.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@41177.4]
  assign RootController_kernelRootController_concrete1_io_in_x202_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 60:23:@41243.4]
  assign RootController_kernelRootController_concrete1_io_in_x201_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 61:23:@41253.4]
  assign RootController_kernelRootController_concrete1_io_in_x201_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 61:23:@41251.4]
  assign RootController_kernelRootController_concrete1_io_in_x201_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 61:23:@41247.4]
  assign RootController_kernelRootController_concrete1_io_in_x201_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 61:23:@41246.4]
  assign RootController_kernelRootController_concrete1_io_in_x361_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 62:23:@41257.4]
  assign RootController_kernelRootController_concrete1_io_in_x360_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 63:23:@41261.4]
  assign RootController_kernelRootController_concrete1_io_in_x362_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 64:23:@41263.4]
  assign RootController_kernelRootController_concrete1_io_in_x199_outdram_number = io_argIns_1; // @[sm_RootController.scala 65:31:@41265.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@41274.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@41272.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@41266.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@41295.2]
  input        clock, // @[:@41296.4]
  input        reset, // @[:@41297.4]
  input        io_enable, // @[:@41298.4]
  output [5:0] io_out, // @[:@41298.4]
  output [5:0] io_next // @[:@41298.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@41300.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@41301.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@41302.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@41307.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@41301.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@41302.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@41307.6]
  assign io_out = count; // @[Counter.scala 25:10:@41310.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@41311.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_25( // @[:@41347.2]
  input         clock, // @[:@41348.4]
  input         reset, // @[:@41349.4]
  input  [5:0]  io_raddr, // @[:@41350.4]
  input         io_wen, // @[:@41350.4]
  input  [5:0]  io_waddr, // @[:@41350.4]
  input  [63:0] io_wdata_addr, // @[:@41350.4]
  input  [31:0] io_wdata_size, // @[:@41350.4]
  output [63:0] io_rdata_addr, // @[:@41350.4]
  output [31:0] io_rdata_size // @[:@41350.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@41352.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@41352.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@41352.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@41352.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@41352.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@41352.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@41352.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@41352.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@41352.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@41366.4]
  wire  _T_20; // @[SRAM.scala 182:49:@41371.4]
  wire  _T_21; // @[SRAM.scala 182:37:@41372.4]
  reg  _T_24; // @[SRAM.scala 182:29:@41373.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@41376.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@41378.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@41352.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@41366.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@41371.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@41372.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@41378.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@41387.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@41386.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@41367.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@41368.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@41364.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@41370.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@41369.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@41365.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@41363.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@41362.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@41389.2]
  input         clock, // @[:@41390.4]
  input         reset, // @[:@41391.4]
  output        io_in_ready, // @[:@41392.4]
  input         io_in_valid, // @[:@41392.4]
  input  [63:0] io_in_bits_addr, // @[:@41392.4]
  input  [31:0] io_in_bits_size, // @[:@41392.4]
  input         io_out_ready, // @[:@41392.4]
  output        io_out_valid, // @[:@41392.4]
  output [63:0] io_out_bits_addr, // @[:@41392.4]
  output [31:0] io_out_bits_size // @[:@41392.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@41788.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@41788.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@41788.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@41788.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@41788.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@41798.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@41798.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@41798.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@41798.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@41798.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@41813.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@41813.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@41813.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@41813.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@41813.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@41813.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@41813.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@41813.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@41813.4]
  wire  writeEn; // @[FIFO.scala 30:29:@41786.4]
  wire  readEn; // @[FIFO.scala 31:29:@41787.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@41808.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@41809.4]
  wire  _T_824; // @[FIFO.scala 45:27:@41810.4]
  wire  empty; // @[FIFO.scala 45:24:@41811.4]
  wire  full; // @[FIFO.scala 46:23:@41812.4]
  wire  _T_827; // @[FIFO.scala 83:17:@41825.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@41826.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@41788.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@41798.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_25 SRAM ( // @[FIFO.scala 73:19:@41813.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@41786.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@41787.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@41809.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@41810.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@41811.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@41812.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@41825.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@41826.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@41832.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@41830.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@41823.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@41822.4]
  assign enqCounter_clock = clock; // @[:@41789.4]
  assign enqCounter_reset = reset; // @[:@41790.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@41796.4]
  assign deqCounter_clock = clock; // @[:@41799.4]
  assign deqCounter_reset = reset; // @[:@41800.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@41806.4]
  assign SRAM_clock = clock; // @[:@41814.4]
  assign SRAM_reset = reset; // @[:@41815.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@41817.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@41818.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@41819.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@41821.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@41820.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@41834.2]
  input        clock, // @[:@41835.4]
  input        reset, // @[:@41836.4]
  input        io_enable, // @[:@41837.4]
  output [3:0] io_out // @[:@41837.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@41839.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@41840.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@41841.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@41846.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@41840.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@41841.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@41846.6]
  assign io_out = count; // @[Counter.scala 25:10:@41849.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@41870.2]
  input        clock, // @[:@41871.4]
  input        reset, // @[:@41872.4]
  input        io_reset, // @[:@41873.4]
  input        io_enable, // @[:@41873.4]
  input  [1:0] io_stride, // @[:@41873.4]
  output [1:0] io_out, // @[:@41873.4]
  output [1:0] io_next // @[:@41873.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@41875.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@41876.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@41877.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@41882.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@41878.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@41876.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@41877.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@41882.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@41878.4]
  assign io_out = count; // @[Counter.scala 25:10:@41885.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@41886.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_26( // @[:@41922.2]
  input         clock, // @[:@41923.4]
  input         reset, // @[:@41924.4]
  input  [1:0]  io_raddr, // @[:@41925.4]
  input         io_wen, // @[:@41925.4]
  input  [1:0]  io_waddr, // @[:@41925.4]
  input  [31:0] io_wdata, // @[:@41925.4]
  output [31:0] io_rdata, // @[:@41925.4]
  input         io_backpressure // @[:@41925.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@41927.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@41927.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@41927.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@41927.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@41927.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@41927.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@41927.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@41927.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@41927.4]
  wire  _T_19; // @[SRAM.scala 182:49:@41945.4]
  wire  _T_20; // @[SRAM.scala 182:37:@41946.4]
  reg  _T_23; // @[SRAM.scala 182:29:@41947.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@41949.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@41927.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@41945.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@41946.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@41954.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@41941.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@41942.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@41939.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@41944.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@41943.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@41940.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@41938.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@41937.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@41956.2]
  input         clock, // @[:@41957.4]
  input         reset, // @[:@41958.4]
  output        io_in_ready, // @[:@41959.4]
  input         io_in_valid, // @[:@41959.4]
  input  [31:0] io_in_bits, // @[:@41959.4]
  input         io_out_ready, // @[:@41959.4]
  output        io_out_valid, // @[:@41959.4]
  output [31:0] io_out_bits // @[:@41959.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@41985.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@41985.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@41985.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@41985.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@41985.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@41985.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@41985.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@41995.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@41995.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@41995.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@41995.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@41995.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@41995.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@41995.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@42010.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@42010.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@42010.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@42010.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@42010.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@42010.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@42010.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@42010.4]
  wire  writeEn; // @[FIFO.scala 30:29:@41983.4]
  wire  readEn; // @[FIFO.scala 31:29:@41984.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@42005.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@42006.4]
  wire  _T_104; // @[FIFO.scala 45:27:@42007.4]
  wire  empty; // @[FIFO.scala 45:24:@42008.4]
  wire  full; // @[FIFO.scala 46:23:@42009.4]
  wire  _T_107; // @[FIFO.scala 83:17:@42020.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@42021.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@41985.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@41995.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_26 SRAM ( // @[FIFO.scala 73:19:@42010.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@41983.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@41984.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@42006.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@42007.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@42008.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@42009.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@42020.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@42021.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@42027.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@42025.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@42018.4]
  assign enqCounter_clock = clock; // @[:@41986.4]
  assign enqCounter_reset = reset; // @[:@41987.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@41993.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@41994.4]
  assign deqCounter_clock = clock; // @[:@41996.4]
  assign deqCounter_reset = reset; // @[:@41997.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@42003.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@42004.4]
  assign SRAM_clock = clock; // @[:@42011.4]
  assign SRAM_reset = reset; // @[:@42012.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@42014.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@42015.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@42016.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@42017.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@42019.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@44414.2]
  input         clock, // @[:@44415.4]
  input         reset, // @[:@44416.4]
  output        io_in_ready, // @[:@44417.4]
  input         io_in_valid, // @[:@44417.4]
  input  [31:0] io_in_bits_0, // @[:@44417.4]
  input         io_out_ready, // @[:@44417.4]
  output        io_out_valid, // @[:@44417.4]
  output [31:0] io_out_bits_0, // @[:@44417.4]
  output [31:0] io_out_bits_1, // @[:@44417.4]
  output [31:0] io_out_bits_2, // @[:@44417.4]
  output [31:0] io_out_bits_3, // @[:@44417.4]
  output [31:0] io_out_bits_4, // @[:@44417.4]
  output [31:0] io_out_bits_5, // @[:@44417.4]
  output [31:0] io_out_bits_6, // @[:@44417.4]
  output [31:0] io_out_bits_7, // @[:@44417.4]
  output [31:0] io_out_bits_8, // @[:@44417.4]
  output [31:0] io_out_bits_9, // @[:@44417.4]
  output [31:0] io_out_bits_10, // @[:@44417.4]
  output [31:0] io_out_bits_11, // @[:@44417.4]
  output [31:0] io_out_bits_12, // @[:@44417.4]
  output [31:0] io_out_bits_13, // @[:@44417.4]
  output [31:0] io_out_bits_14, // @[:@44417.4]
  output [31:0] io_out_bits_15 // @[:@44417.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@44421.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@44421.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@44421.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@44421.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@44432.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@44432.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@44432.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@44432.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@44445.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@44445.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@44445.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@44445.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@44445.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@44445.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@44445.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@44445.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@44480.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@44480.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@44480.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@44480.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@44480.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@44480.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@44480.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@44480.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@44515.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@44515.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@44515.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@44515.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@44515.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@44515.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@44515.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@44515.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@44550.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@44550.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@44550.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@44550.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@44550.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@44550.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@44550.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@44550.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@44585.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@44585.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@44585.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@44585.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@44585.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@44585.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@44585.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@44585.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@44620.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@44620.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@44620.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@44620.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@44620.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@44620.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@44620.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@44620.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@44655.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@44655.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@44655.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@44655.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@44655.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@44655.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@44655.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@44655.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@44690.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@44690.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@44690.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@44690.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@44690.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@44690.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@44690.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@44690.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@44725.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@44725.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@44725.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@44725.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@44725.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@44725.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@44725.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@44725.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@44760.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@44760.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@44760.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@44760.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@44760.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@44760.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@44760.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@44760.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@44795.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@44795.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@44795.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@44795.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@44795.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@44795.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@44795.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@44795.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@44830.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@44830.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@44830.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@44830.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@44830.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@44830.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@44830.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@44830.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@44865.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@44865.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@44865.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@44865.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@44865.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@44865.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@44865.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@44865.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@44900.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@44900.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@44900.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@44900.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@44900.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@44900.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@44900.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@44900.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@44935.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@44935.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@44935.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@44935.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@44935.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@44935.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@44935.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@44935.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@44970.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@44970.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@44970.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@44970.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@44970.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@44970.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@44970.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@44970.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@44420.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@44443.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@44470.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@44505.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@44540.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@44575.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@44610.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@44645.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@44680.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@44715.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@44750.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@44785.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@44820.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@44855.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@44890.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@44925.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@44960.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@44995.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45006.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45007.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45008.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45009.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45010.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45011.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45012.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45013.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45014.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45015.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45016.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45017.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45018.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45019.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45020.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@45037.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45021.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@45056.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@45057.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@45058.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@45059.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@45060.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@45061.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@45062.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@45063.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@45064.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@45065.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@45066.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@45067.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@45068.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@45069.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@44421.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@44432.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@44445.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@44480.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@44515.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@44550.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@44585.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@44620.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@44655.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@44690.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@44725.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@44760.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@44795.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@44830.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@44865.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@44900.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@44935.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@44970.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@44420.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@44443.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@44470.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@44505.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@44540.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@44575.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@44610.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@44645.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@44680.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@44715.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@44750.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@44785.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@44820.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@44855.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@44890.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@44925.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@44960.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@44995.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45006.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45007.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45008.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45009.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45010.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45011.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45012.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45013.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45014.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45015.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45016.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45017.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45018.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45019.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45020.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@45037.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@45005.4 FIFOVec.scala 49:42:@45021.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@45056.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@45057.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@45058.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@45059.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@45060.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@45061.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@45062.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@45063.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@45064.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@45065.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@45066.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@45067.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@45068.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@45069.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@45038.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@45072.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@45380.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@45381.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@45382.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@45383.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@45384.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@45385.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@45386.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@45387.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@45388.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@45389.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@45390.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@45391.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@45392.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@45393.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@45394.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@45395.4]
  assign enqCounter_clock = clock; // @[:@44422.4]
  assign enqCounter_reset = reset; // @[:@44423.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@44430.4]
  assign deqCounter_clock = clock; // @[:@44433.4]
  assign deqCounter_reset = reset; // @[:@44434.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@44441.4]
  assign fifos_0_clock = clock; // @[:@44446.4]
  assign fifos_0_reset = reset; // @[:@44447.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@44473.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44475.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44479.4]
  assign fifos_1_clock = clock; // @[:@44481.4]
  assign fifos_1_reset = reset; // @[:@44482.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@44508.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44510.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44514.4]
  assign fifos_2_clock = clock; // @[:@44516.4]
  assign fifos_2_reset = reset; // @[:@44517.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@44543.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44545.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44549.4]
  assign fifos_3_clock = clock; // @[:@44551.4]
  assign fifos_3_reset = reset; // @[:@44552.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@44578.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44580.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44584.4]
  assign fifos_4_clock = clock; // @[:@44586.4]
  assign fifos_4_reset = reset; // @[:@44587.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@44613.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44615.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44619.4]
  assign fifos_5_clock = clock; // @[:@44621.4]
  assign fifos_5_reset = reset; // @[:@44622.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@44648.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44650.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44654.4]
  assign fifos_6_clock = clock; // @[:@44656.4]
  assign fifos_6_reset = reset; // @[:@44657.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@44683.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44685.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44689.4]
  assign fifos_7_clock = clock; // @[:@44691.4]
  assign fifos_7_reset = reset; // @[:@44692.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@44718.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44720.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44724.4]
  assign fifos_8_clock = clock; // @[:@44726.4]
  assign fifos_8_reset = reset; // @[:@44727.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@44753.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44755.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44759.4]
  assign fifos_9_clock = clock; // @[:@44761.4]
  assign fifos_9_reset = reset; // @[:@44762.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@44788.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44790.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44794.4]
  assign fifos_10_clock = clock; // @[:@44796.4]
  assign fifos_10_reset = reset; // @[:@44797.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@44823.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44825.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44829.4]
  assign fifos_11_clock = clock; // @[:@44831.4]
  assign fifos_11_reset = reset; // @[:@44832.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@44858.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44860.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44864.4]
  assign fifos_12_clock = clock; // @[:@44866.4]
  assign fifos_12_reset = reset; // @[:@44867.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@44893.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44895.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44899.4]
  assign fifos_13_clock = clock; // @[:@44901.4]
  assign fifos_13_reset = reset; // @[:@44902.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@44928.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44930.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44934.4]
  assign fifos_14_clock = clock; // @[:@44936.4]
  assign fifos_14_reset = reset; // @[:@44937.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@44963.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44965.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44969.4]
  assign fifos_15_clock = clock; // @[:@44971.4]
  assign fifos_15_reset = reset; // @[:@44972.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@44998.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@45000.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@45004.4]
endmodule
module FFRAM( // @[:@45469.2]
  input        clock, // @[:@45470.4]
  input        reset, // @[:@45471.4]
  input  [1:0] io_raddr, // @[:@45472.4]
  input        io_wen, // @[:@45472.4]
  input  [1:0] io_waddr, // @[:@45472.4]
  input        io_wdata, // @[:@45472.4]
  output       io_rdata, // @[:@45472.4]
  input        io_banks_0_wdata_valid, // @[:@45472.4]
  input        io_banks_0_wdata_bits, // @[:@45472.4]
  input        io_banks_1_wdata_valid, // @[:@45472.4]
  input        io_banks_1_wdata_bits, // @[:@45472.4]
  input        io_banks_2_wdata_valid, // @[:@45472.4]
  input        io_banks_2_wdata_bits, // @[:@45472.4]
  input        io_banks_3_wdata_valid, // @[:@45472.4]
  input        io_banks_3_wdata_bits // @[:@45472.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@45476.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@45477.4]
  wire  _T_89; // @[SRAM.scala 148:25:@45478.4]
  wire  _T_90; // @[SRAM.scala 148:15:@45479.4]
  wire  _T_91; // @[SRAM.scala 149:15:@45481.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@45480.4]
  reg  regs_1; // @[SRAM.scala 145:20:@45487.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@45488.4]
  wire  _T_98; // @[SRAM.scala 148:25:@45489.4]
  wire  _T_99; // @[SRAM.scala 148:15:@45490.4]
  wire  _T_100; // @[SRAM.scala 149:15:@45492.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@45491.4]
  reg  regs_2; // @[SRAM.scala 145:20:@45498.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@45499.4]
  wire  _T_107; // @[SRAM.scala 148:25:@45500.4]
  wire  _T_108; // @[SRAM.scala 148:15:@45501.4]
  wire  _T_109; // @[SRAM.scala 149:15:@45503.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@45502.4]
  reg  regs_3; // @[SRAM.scala 145:20:@45509.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@45510.4]
  wire  _T_116; // @[SRAM.scala 148:25:@45511.4]
  wire  _T_117; // @[SRAM.scala 148:15:@45512.4]
  wire  _T_118; // @[SRAM.scala 149:15:@45514.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@45513.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@45523.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@45523.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@45477.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@45478.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@45479.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45481.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@45480.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@45488.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@45489.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@45490.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45492.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@45491.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@45499.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@45500.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@45501.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45503.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@45502.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@45510.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@45511.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@45512.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45514.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@45513.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@45523.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@45523.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@45523.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@45525.2]
  input   clock, // @[:@45526.4]
  input   reset, // @[:@45527.4]
  output  io_in_ready, // @[:@45528.4]
  input   io_in_valid, // @[:@45528.4]
  input   io_in_bits, // @[:@45528.4]
  input   io_out_ready, // @[:@45528.4]
  output  io_out_valid, // @[:@45528.4]
  output  io_out_bits // @[:@45528.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@45554.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@45554.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@45554.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@45554.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@45554.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@45554.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@45554.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@45564.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@45564.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@45564.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@45564.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@45564.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@45564.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@45564.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@45579.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@45579.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@45579.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@45579.4]
  wire  writeEn; // @[FIFO.scala 30:29:@45552.4]
  wire  readEn; // @[FIFO.scala 31:29:@45553.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@45574.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@45575.4]
  wire  _T_104; // @[FIFO.scala 45:27:@45576.4]
  wire  empty; // @[FIFO.scala 45:24:@45577.4]
  wire  full; // @[FIFO.scala 46:23:@45578.4]
  wire  _T_157; // @[FIFO.scala 83:17:@45665.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@45666.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@45554.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@45564.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@45579.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@45552.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@45553.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@45575.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@45576.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@45577.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@45578.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@45665.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@45666.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@45672.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@45670.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@45604.4]
  assign enqCounter_clock = clock; // @[:@45555.4]
  assign enqCounter_reset = reset; // @[:@45556.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@45562.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@45563.4]
  assign deqCounter_clock = clock; // @[:@45565.4]
  assign deqCounter_reset = reset; // @[:@45566.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@45572.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@45573.4]
  assign FFRAM_clock = clock; // @[:@45580.4]
  assign FFRAM_reset = reset; // @[:@45581.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@45600.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@45601.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@45602.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@45603.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45606.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45605.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45609.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45608.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45612.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45611.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45615.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45614.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@49289.2]
  input   clock, // @[:@49290.4]
  input   reset, // @[:@49291.4]
  output  io_in_ready, // @[:@49292.4]
  input   io_in_valid, // @[:@49292.4]
  input   io_in_bits_0, // @[:@49292.4]
  input   io_out_ready, // @[:@49292.4]
  output  io_out_valid, // @[:@49292.4]
  output  io_out_bits_0, // @[:@49292.4]
  output  io_out_bits_1, // @[:@49292.4]
  output  io_out_bits_2, // @[:@49292.4]
  output  io_out_bits_3, // @[:@49292.4]
  output  io_out_bits_4, // @[:@49292.4]
  output  io_out_bits_5, // @[:@49292.4]
  output  io_out_bits_6, // @[:@49292.4]
  output  io_out_bits_7, // @[:@49292.4]
  output  io_out_bits_8, // @[:@49292.4]
  output  io_out_bits_9, // @[:@49292.4]
  output  io_out_bits_10, // @[:@49292.4]
  output  io_out_bits_11, // @[:@49292.4]
  output  io_out_bits_12, // @[:@49292.4]
  output  io_out_bits_13, // @[:@49292.4]
  output  io_out_bits_14, // @[:@49292.4]
  output  io_out_bits_15 // @[:@49292.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@49296.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@49296.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@49296.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@49296.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@49307.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@49307.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@49307.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@49307.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@49320.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@49355.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@49390.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@49425.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@49460.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@49495.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@49530.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@49565.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@49600.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@49635.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@49670.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@49705.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@49740.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@49775.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@49810.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@49845.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@49845.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@49845.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@49845.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@49845.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@49845.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@49845.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@49845.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@49295.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@49318.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@49345.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@49380.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@49415.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@49450.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@49485.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@49520.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@49555.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@49590.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@49625.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@49660.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@49695.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@49730.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@49765.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@49800.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@49835.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@49870.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49881.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49882.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49883.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49884.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49885.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49886.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49887.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49888.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49889.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49890.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49891.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49892.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49893.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49894.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49895.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@49912.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49896.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@49931.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@49932.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@49933.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@49934.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@49935.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@49936.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@49937.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@49938.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@49939.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@49940.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@49941.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@49942.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@49943.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@49944.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@49296.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@49307.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@49320.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@49355.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@49390.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@49425.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@49460.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@49495.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@49530.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@49565.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@49600.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@49635.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@49670.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@49705.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@49740.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@49775.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@49810.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@49845.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@49295.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@49318.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@49345.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@49380.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@49415.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@49450.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@49485.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@49520.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@49555.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@49590.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@49625.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@49660.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@49695.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@49730.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@49765.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@49800.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@49835.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@49870.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49881.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49882.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49883.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49884.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49885.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49886.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49887.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49888.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49889.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49890.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49891.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49892.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49893.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49894.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49895.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@49912.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@49880.4 FIFOVec.scala 49:42:@49896.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@49931.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@49932.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@49933.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@49934.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@49935.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@49936.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@49937.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@49938.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@49939.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@49940.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@49941.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@49942.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@49943.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@49944.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@49913.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@49947.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@50255.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@50256.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@50257.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@50258.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@50259.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@50260.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@50261.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@50262.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@50263.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@50264.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@50265.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@50266.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@50267.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@50268.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@50269.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@50270.4]
  assign enqCounter_clock = clock; // @[:@49297.4]
  assign enqCounter_reset = reset; // @[:@49298.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@49305.4]
  assign deqCounter_clock = clock; // @[:@49308.4]
  assign deqCounter_reset = reset; // @[:@49309.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@49316.4]
  assign fifos_0_clock = clock; // @[:@49321.4]
  assign fifos_0_reset = reset; // @[:@49322.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@49348.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49350.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49354.4]
  assign fifos_1_clock = clock; // @[:@49356.4]
  assign fifos_1_reset = reset; // @[:@49357.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@49383.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49385.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49389.4]
  assign fifos_2_clock = clock; // @[:@49391.4]
  assign fifos_2_reset = reset; // @[:@49392.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@49418.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49420.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49424.4]
  assign fifos_3_clock = clock; // @[:@49426.4]
  assign fifos_3_reset = reset; // @[:@49427.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@49453.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49455.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49459.4]
  assign fifos_4_clock = clock; // @[:@49461.4]
  assign fifos_4_reset = reset; // @[:@49462.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@49488.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49490.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49494.4]
  assign fifos_5_clock = clock; // @[:@49496.4]
  assign fifos_5_reset = reset; // @[:@49497.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@49523.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49525.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49529.4]
  assign fifos_6_clock = clock; // @[:@49531.4]
  assign fifos_6_reset = reset; // @[:@49532.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@49558.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49560.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49564.4]
  assign fifos_7_clock = clock; // @[:@49566.4]
  assign fifos_7_reset = reset; // @[:@49567.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@49593.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49595.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49599.4]
  assign fifos_8_clock = clock; // @[:@49601.4]
  assign fifos_8_reset = reset; // @[:@49602.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@49628.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49630.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49634.4]
  assign fifos_9_clock = clock; // @[:@49636.4]
  assign fifos_9_reset = reset; // @[:@49637.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@49663.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49665.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49669.4]
  assign fifos_10_clock = clock; // @[:@49671.4]
  assign fifos_10_reset = reset; // @[:@49672.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@49698.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49700.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49704.4]
  assign fifos_11_clock = clock; // @[:@49706.4]
  assign fifos_11_reset = reset; // @[:@49707.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@49733.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49735.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49739.4]
  assign fifos_12_clock = clock; // @[:@49741.4]
  assign fifos_12_reset = reset; // @[:@49742.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@49768.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49770.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49774.4]
  assign fifos_13_clock = clock; // @[:@49776.4]
  assign fifos_13_reset = reset; // @[:@49777.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@49803.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49805.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49809.4]
  assign fifos_14_clock = clock; // @[:@49811.4]
  assign fifos_14_reset = reset; // @[:@49812.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@49838.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49840.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49844.4]
  assign fifos_15_clock = clock; // @[:@49846.4]
  assign fifos_15_reset = reset; // @[:@49847.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@49873.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49875.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49879.4]
endmodule
module FIFOWidthConvert( // @[:@50272.2]
  input         clock, // @[:@50273.4]
  input         reset, // @[:@50274.4]
  output        io_in_ready, // @[:@50275.4]
  input         io_in_valid, // @[:@50275.4]
  input  [31:0] io_in_bits_data_0, // @[:@50275.4]
  input         io_in_bits_strobe, // @[:@50275.4]
  input         io_out_ready, // @[:@50275.4]
  output        io_out_valid, // @[:@50275.4]
  output [31:0] io_out_bits_data_0, // @[:@50275.4]
  output [31:0] io_out_bits_data_1, // @[:@50275.4]
  output [31:0] io_out_bits_data_2, // @[:@50275.4]
  output [31:0] io_out_bits_data_3, // @[:@50275.4]
  output [31:0] io_out_bits_data_4, // @[:@50275.4]
  output [31:0] io_out_bits_data_5, // @[:@50275.4]
  output [31:0] io_out_bits_data_6, // @[:@50275.4]
  output [31:0] io_out_bits_data_7, // @[:@50275.4]
  output [31:0] io_out_bits_data_8, // @[:@50275.4]
  output [31:0] io_out_bits_data_9, // @[:@50275.4]
  output [31:0] io_out_bits_data_10, // @[:@50275.4]
  output [31:0] io_out_bits_data_11, // @[:@50275.4]
  output [31:0] io_out_bits_data_12, // @[:@50275.4]
  output [31:0] io_out_bits_data_13, // @[:@50275.4]
  output [31:0] io_out_bits_data_14, // @[:@50275.4]
  output [31:0] io_out_bits_data_15, // @[:@50275.4]
  output [63:0] io_out_bits_strobe // @[:@50275.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@50277.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@50318.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@50377.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@50383.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@50441.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@50447.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@50448.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@50452.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@50456.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@50460.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@50464.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@50468.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@50472.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@50476.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@50480.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@50484.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@50488.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@50492.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@50496.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@50500.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@50504.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@50508.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@50585.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@50594.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@50603.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@50612.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@50621.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@50630.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@50638.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@50277.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@50318.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@50377.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@50383.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@50441.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@50447.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@50448.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@50452.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@50456.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@50460.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@50464.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@50468.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@50472.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@50476.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@50480.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@50484.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@50488.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@50492.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@50496.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@50500.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@50504.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@50508.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@50585.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@50594.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@50603.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@50612.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@50621.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@50630.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@50638.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@50367.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@50368.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@50417.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@50418.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@50419.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@50420.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@50421.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@50422.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@50423.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@50424.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@50425.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@50426.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@50427.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@50428.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@50429.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@50430.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@50431.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@50432.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@50640.4]
  assign FIFOVec_clock = clock; // @[:@50278.4]
  assign FIFOVec_reset = reset; // @[:@50279.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@50364.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@50363.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@50641.4]
  assign FIFOVec_1_clock = clock; // @[:@50319.4]
  assign FIFOVec_1_reset = reset; // @[:@50320.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@50366.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@50365.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@50642.4]
endmodule
module FFRAM_16( // @[:@50680.2]
  input        clock, // @[:@50681.4]
  input        reset, // @[:@50682.4]
  input  [5:0] io_raddr, // @[:@50683.4]
  input        io_wen, // @[:@50683.4]
  input  [5:0] io_waddr, // @[:@50683.4]
  input        io_wdata, // @[:@50683.4]
  output       io_rdata, // @[:@50683.4]
  input        io_banks_0_wdata_valid, // @[:@50683.4]
  input        io_banks_0_wdata_bits, // @[:@50683.4]
  input        io_banks_1_wdata_valid, // @[:@50683.4]
  input        io_banks_1_wdata_bits, // @[:@50683.4]
  input        io_banks_2_wdata_valid, // @[:@50683.4]
  input        io_banks_2_wdata_bits, // @[:@50683.4]
  input        io_banks_3_wdata_valid, // @[:@50683.4]
  input        io_banks_3_wdata_bits, // @[:@50683.4]
  input        io_banks_4_wdata_valid, // @[:@50683.4]
  input        io_banks_4_wdata_bits, // @[:@50683.4]
  input        io_banks_5_wdata_valid, // @[:@50683.4]
  input        io_banks_5_wdata_bits, // @[:@50683.4]
  input        io_banks_6_wdata_valid, // @[:@50683.4]
  input        io_banks_6_wdata_bits, // @[:@50683.4]
  input        io_banks_7_wdata_valid, // @[:@50683.4]
  input        io_banks_7_wdata_bits, // @[:@50683.4]
  input        io_banks_8_wdata_valid, // @[:@50683.4]
  input        io_banks_8_wdata_bits, // @[:@50683.4]
  input        io_banks_9_wdata_valid, // @[:@50683.4]
  input        io_banks_9_wdata_bits, // @[:@50683.4]
  input        io_banks_10_wdata_valid, // @[:@50683.4]
  input        io_banks_10_wdata_bits, // @[:@50683.4]
  input        io_banks_11_wdata_valid, // @[:@50683.4]
  input        io_banks_11_wdata_bits, // @[:@50683.4]
  input        io_banks_12_wdata_valid, // @[:@50683.4]
  input        io_banks_12_wdata_bits, // @[:@50683.4]
  input        io_banks_13_wdata_valid, // @[:@50683.4]
  input        io_banks_13_wdata_bits, // @[:@50683.4]
  input        io_banks_14_wdata_valid, // @[:@50683.4]
  input        io_banks_14_wdata_bits, // @[:@50683.4]
  input        io_banks_15_wdata_valid, // @[:@50683.4]
  input        io_banks_15_wdata_bits, // @[:@50683.4]
  input        io_banks_16_wdata_valid, // @[:@50683.4]
  input        io_banks_16_wdata_bits, // @[:@50683.4]
  input        io_banks_17_wdata_valid, // @[:@50683.4]
  input        io_banks_17_wdata_bits, // @[:@50683.4]
  input        io_banks_18_wdata_valid, // @[:@50683.4]
  input        io_banks_18_wdata_bits, // @[:@50683.4]
  input        io_banks_19_wdata_valid, // @[:@50683.4]
  input        io_banks_19_wdata_bits, // @[:@50683.4]
  input        io_banks_20_wdata_valid, // @[:@50683.4]
  input        io_banks_20_wdata_bits, // @[:@50683.4]
  input        io_banks_21_wdata_valid, // @[:@50683.4]
  input        io_banks_21_wdata_bits, // @[:@50683.4]
  input        io_banks_22_wdata_valid, // @[:@50683.4]
  input        io_banks_22_wdata_bits, // @[:@50683.4]
  input        io_banks_23_wdata_valid, // @[:@50683.4]
  input        io_banks_23_wdata_bits, // @[:@50683.4]
  input        io_banks_24_wdata_valid, // @[:@50683.4]
  input        io_banks_24_wdata_bits, // @[:@50683.4]
  input        io_banks_25_wdata_valid, // @[:@50683.4]
  input        io_banks_25_wdata_bits, // @[:@50683.4]
  input        io_banks_26_wdata_valid, // @[:@50683.4]
  input        io_banks_26_wdata_bits, // @[:@50683.4]
  input        io_banks_27_wdata_valid, // @[:@50683.4]
  input        io_banks_27_wdata_bits, // @[:@50683.4]
  input        io_banks_28_wdata_valid, // @[:@50683.4]
  input        io_banks_28_wdata_bits, // @[:@50683.4]
  input        io_banks_29_wdata_valid, // @[:@50683.4]
  input        io_banks_29_wdata_bits, // @[:@50683.4]
  input        io_banks_30_wdata_valid, // @[:@50683.4]
  input        io_banks_30_wdata_bits, // @[:@50683.4]
  input        io_banks_31_wdata_valid, // @[:@50683.4]
  input        io_banks_31_wdata_bits, // @[:@50683.4]
  input        io_banks_32_wdata_valid, // @[:@50683.4]
  input        io_banks_32_wdata_bits, // @[:@50683.4]
  input        io_banks_33_wdata_valid, // @[:@50683.4]
  input        io_banks_33_wdata_bits, // @[:@50683.4]
  input        io_banks_34_wdata_valid, // @[:@50683.4]
  input        io_banks_34_wdata_bits, // @[:@50683.4]
  input        io_banks_35_wdata_valid, // @[:@50683.4]
  input        io_banks_35_wdata_bits, // @[:@50683.4]
  input        io_banks_36_wdata_valid, // @[:@50683.4]
  input        io_banks_36_wdata_bits, // @[:@50683.4]
  input        io_banks_37_wdata_valid, // @[:@50683.4]
  input        io_banks_37_wdata_bits, // @[:@50683.4]
  input        io_banks_38_wdata_valid, // @[:@50683.4]
  input        io_banks_38_wdata_bits, // @[:@50683.4]
  input        io_banks_39_wdata_valid, // @[:@50683.4]
  input        io_banks_39_wdata_bits, // @[:@50683.4]
  input        io_banks_40_wdata_valid, // @[:@50683.4]
  input        io_banks_40_wdata_bits, // @[:@50683.4]
  input        io_banks_41_wdata_valid, // @[:@50683.4]
  input        io_banks_41_wdata_bits, // @[:@50683.4]
  input        io_banks_42_wdata_valid, // @[:@50683.4]
  input        io_banks_42_wdata_bits, // @[:@50683.4]
  input        io_banks_43_wdata_valid, // @[:@50683.4]
  input        io_banks_43_wdata_bits, // @[:@50683.4]
  input        io_banks_44_wdata_valid, // @[:@50683.4]
  input        io_banks_44_wdata_bits, // @[:@50683.4]
  input        io_banks_45_wdata_valid, // @[:@50683.4]
  input        io_banks_45_wdata_bits, // @[:@50683.4]
  input        io_banks_46_wdata_valid, // @[:@50683.4]
  input        io_banks_46_wdata_bits, // @[:@50683.4]
  input        io_banks_47_wdata_valid, // @[:@50683.4]
  input        io_banks_47_wdata_bits, // @[:@50683.4]
  input        io_banks_48_wdata_valid, // @[:@50683.4]
  input        io_banks_48_wdata_bits, // @[:@50683.4]
  input        io_banks_49_wdata_valid, // @[:@50683.4]
  input        io_banks_49_wdata_bits, // @[:@50683.4]
  input        io_banks_50_wdata_valid, // @[:@50683.4]
  input        io_banks_50_wdata_bits, // @[:@50683.4]
  input        io_banks_51_wdata_valid, // @[:@50683.4]
  input        io_banks_51_wdata_bits, // @[:@50683.4]
  input        io_banks_52_wdata_valid, // @[:@50683.4]
  input        io_banks_52_wdata_bits, // @[:@50683.4]
  input        io_banks_53_wdata_valid, // @[:@50683.4]
  input        io_banks_53_wdata_bits, // @[:@50683.4]
  input        io_banks_54_wdata_valid, // @[:@50683.4]
  input        io_banks_54_wdata_bits, // @[:@50683.4]
  input        io_banks_55_wdata_valid, // @[:@50683.4]
  input        io_banks_55_wdata_bits, // @[:@50683.4]
  input        io_banks_56_wdata_valid, // @[:@50683.4]
  input        io_banks_56_wdata_bits, // @[:@50683.4]
  input        io_banks_57_wdata_valid, // @[:@50683.4]
  input        io_banks_57_wdata_bits, // @[:@50683.4]
  input        io_banks_58_wdata_valid, // @[:@50683.4]
  input        io_banks_58_wdata_bits, // @[:@50683.4]
  input        io_banks_59_wdata_valid, // @[:@50683.4]
  input        io_banks_59_wdata_bits, // @[:@50683.4]
  input        io_banks_60_wdata_valid, // @[:@50683.4]
  input        io_banks_60_wdata_bits, // @[:@50683.4]
  input        io_banks_61_wdata_valid, // @[:@50683.4]
  input        io_banks_61_wdata_bits, // @[:@50683.4]
  input        io_banks_62_wdata_valid, // @[:@50683.4]
  input        io_banks_62_wdata_bits, // @[:@50683.4]
  input        io_banks_63_wdata_valid, // @[:@50683.4]
  input        io_banks_63_wdata_bits // @[:@50683.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@50687.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@50688.4]
  wire  _T_689; // @[SRAM.scala 148:25:@50689.4]
  wire  _T_690; // @[SRAM.scala 148:15:@50690.4]
  wire  _T_691; // @[SRAM.scala 149:15:@50692.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@50691.4]
  reg  regs_1; // @[SRAM.scala 145:20:@50698.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@50699.4]
  wire  _T_698; // @[SRAM.scala 148:25:@50700.4]
  wire  _T_699; // @[SRAM.scala 148:15:@50701.4]
  wire  _T_700; // @[SRAM.scala 149:15:@50703.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@50702.4]
  reg  regs_2; // @[SRAM.scala 145:20:@50709.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@50710.4]
  wire  _T_707; // @[SRAM.scala 148:25:@50711.4]
  wire  _T_708; // @[SRAM.scala 148:15:@50712.4]
  wire  _T_709; // @[SRAM.scala 149:15:@50714.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@50713.4]
  reg  regs_3; // @[SRAM.scala 145:20:@50720.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@50721.4]
  wire  _T_716; // @[SRAM.scala 148:25:@50722.4]
  wire  _T_717; // @[SRAM.scala 148:15:@50723.4]
  wire  _T_718; // @[SRAM.scala 149:15:@50725.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@50724.4]
  reg  regs_4; // @[SRAM.scala 145:20:@50731.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@50732.4]
  wire  _T_725; // @[SRAM.scala 148:25:@50733.4]
  wire  _T_726; // @[SRAM.scala 148:15:@50734.4]
  wire  _T_727; // @[SRAM.scala 149:15:@50736.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@50735.4]
  reg  regs_5; // @[SRAM.scala 145:20:@50742.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@50743.4]
  wire  _T_734; // @[SRAM.scala 148:25:@50744.4]
  wire  _T_735; // @[SRAM.scala 148:15:@50745.4]
  wire  _T_736; // @[SRAM.scala 149:15:@50747.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@50746.4]
  reg  regs_6; // @[SRAM.scala 145:20:@50753.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@50754.4]
  wire  _T_743; // @[SRAM.scala 148:25:@50755.4]
  wire  _T_744; // @[SRAM.scala 148:15:@50756.4]
  wire  _T_745; // @[SRAM.scala 149:15:@50758.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@50757.4]
  reg  regs_7; // @[SRAM.scala 145:20:@50764.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@50765.4]
  wire  _T_752; // @[SRAM.scala 148:25:@50766.4]
  wire  _T_753; // @[SRAM.scala 148:15:@50767.4]
  wire  _T_754; // @[SRAM.scala 149:15:@50769.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@50768.4]
  reg  regs_8; // @[SRAM.scala 145:20:@50775.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@50776.4]
  wire  _T_761; // @[SRAM.scala 148:25:@50777.4]
  wire  _T_762; // @[SRAM.scala 148:15:@50778.4]
  wire  _T_763; // @[SRAM.scala 149:15:@50780.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@50779.4]
  reg  regs_9; // @[SRAM.scala 145:20:@50786.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@50787.4]
  wire  _T_770; // @[SRAM.scala 148:25:@50788.4]
  wire  _T_771; // @[SRAM.scala 148:15:@50789.4]
  wire  _T_772; // @[SRAM.scala 149:15:@50791.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@50790.4]
  reg  regs_10; // @[SRAM.scala 145:20:@50797.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@50798.4]
  wire  _T_779; // @[SRAM.scala 148:25:@50799.4]
  wire  _T_780; // @[SRAM.scala 148:15:@50800.4]
  wire  _T_781; // @[SRAM.scala 149:15:@50802.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@50801.4]
  reg  regs_11; // @[SRAM.scala 145:20:@50808.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@50809.4]
  wire  _T_788; // @[SRAM.scala 148:25:@50810.4]
  wire  _T_789; // @[SRAM.scala 148:15:@50811.4]
  wire  _T_790; // @[SRAM.scala 149:15:@50813.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@50812.4]
  reg  regs_12; // @[SRAM.scala 145:20:@50819.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@50820.4]
  wire  _T_797; // @[SRAM.scala 148:25:@50821.4]
  wire  _T_798; // @[SRAM.scala 148:15:@50822.4]
  wire  _T_799; // @[SRAM.scala 149:15:@50824.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@50823.4]
  reg  regs_13; // @[SRAM.scala 145:20:@50830.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@50831.4]
  wire  _T_806; // @[SRAM.scala 148:25:@50832.4]
  wire  _T_807; // @[SRAM.scala 148:15:@50833.4]
  wire  _T_808; // @[SRAM.scala 149:15:@50835.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@50834.4]
  reg  regs_14; // @[SRAM.scala 145:20:@50841.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@50842.4]
  wire  _T_815; // @[SRAM.scala 148:25:@50843.4]
  wire  _T_816; // @[SRAM.scala 148:15:@50844.4]
  wire  _T_817; // @[SRAM.scala 149:15:@50846.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@50845.4]
  reg  regs_15; // @[SRAM.scala 145:20:@50852.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@50853.4]
  wire  _T_824; // @[SRAM.scala 148:25:@50854.4]
  wire  _T_825; // @[SRAM.scala 148:15:@50855.4]
  wire  _T_826; // @[SRAM.scala 149:15:@50857.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@50856.4]
  reg  regs_16; // @[SRAM.scala 145:20:@50863.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@50864.4]
  wire  _T_833; // @[SRAM.scala 148:25:@50865.4]
  wire  _T_834; // @[SRAM.scala 148:15:@50866.4]
  wire  _T_835; // @[SRAM.scala 149:15:@50868.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@50867.4]
  reg  regs_17; // @[SRAM.scala 145:20:@50874.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@50875.4]
  wire  _T_842; // @[SRAM.scala 148:25:@50876.4]
  wire  _T_843; // @[SRAM.scala 148:15:@50877.4]
  wire  _T_844; // @[SRAM.scala 149:15:@50879.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@50878.4]
  reg  regs_18; // @[SRAM.scala 145:20:@50885.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@50886.4]
  wire  _T_851; // @[SRAM.scala 148:25:@50887.4]
  wire  _T_852; // @[SRAM.scala 148:15:@50888.4]
  wire  _T_853; // @[SRAM.scala 149:15:@50890.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@50889.4]
  reg  regs_19; // @[SRAM.scala 145:20:@50896.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@50897.4]
  wire  _T_860; // @[SRAM.scala 148:25:@50898.4]
  wire  _T_861; // @[SRAM.scala 148:15:@50899.4]
  wire  _T_862; // @[SRAM.scala 149:15:@50901.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@50900.4]
  reg  regs_20; // @[SRAM.scala 145:20:@50907.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@50908.4]
  wire  _T_869; // @[SRAM.scala 148:25:@50909.4]
  wire  _T_870; // @[SRAM.scala 148:15:@50910.4]
  wire  _T_871; // @[SRAM.scala 149:15:@50912.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@50911.4]
  reg  regs_21; // @[SRAM.scala 145:20:@50918.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@50919.4]
  wire  _T_878; // @[SRAM.scala 148:25:@50920.4]
  wire  _T_879; // @[SRAM.scala 148:15:@50921.4]
  wire  _T_880; // @[SRAM.scala 149:15:@50923.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@50922.4]
  reg  regs_22; // @[SRAM.scala 145:20:@50929.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@50930.4]
  wire  _T_887; // @[SRAM.scala 148:25:@50931.4]
  wire  _T_888; // @[SRAM.scala 148:15:@50932.4]
  wire  _T_889; // @[SRAM.scala 149:15:@50934.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@50933.4]
  reg  regs_23; // @[SRAM.scala 145:20:@50940.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@50941.4]
  wire  _T_896; // @[SRAM.scala 148:25:@50942.4]
  wire  _T_897; // @[SRAM.scala 148:15:@50943.4]
  wire  _T_898; // @[SRAM.scala 149:15:@50945.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@50944.4]
  reg  regs_24; // @[SRAM.scala 145:20:@50951.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@50952.4]
  wire  _T_905; // @[SRAM.scala 148:25:@50953.4]
  wire  _T_906; // @[SRAM.scala 148:15:@50954.4]
  wire  _T_907; // @[SRAM.scala 149:15:@50956.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@50955.4]
  reg  regs_25; // @[SRAM.scala 145:20:@50962.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@50963.4]
  wire  _T_914; // @[SRAM.scala 148:25:@50964.4]
  wire  _T_915; // @[SRAM.scala 148:15:@50965.4]
  wire  _T_916; // @[SRAM.scala 149:15:@50967.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@50966.4]
  reg  regs_26; // @[SRAM.scala 145:20:@50973.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@50974.4]
  wire  _T_923; // @[SRAM.scala 148:25:@50975.4]
  wire  _T_924; // @[SRAM.scala 148:15:@50976.4]
  wire  _T_925; // @[SRAM.scala 149:15:@50978.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@50977.4]
  reg  regs_27; // @[SRAM.scala 145:20:@50984.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@50985.4]
  wire  _T_932; // @[SRAM.scala 148:25:@50986.4]
  wire  _T_933; // @[SRAM.scala 148:15:@50987.4]
  wire  _T_934; // @[SRAM.scala 149:15:@50989.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@50988.4]
  reg  regs_28; // @[SRAM.scala 145:20:@50995.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@50996.4]
  wire  _T_941; // @[SRAM.scala 148:25:@50997.4]
  wire  _T_942; // @[SRAM.scala 148:15:@50998.4]
  wire  _T_943; // @[SRAM.scala 149:15:@51000.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@50999.4]
  reg  regs_29; // @[SRAM.scala 145:20:@51006.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@51007.4]
  wire  _T_950; // @[SRAM.scala 148:25:@51008.4]
  wire  _T_951; // @[SRAM.scala 148:15:@51009.4]
  wire  _T_952; // @[SRAM.scala 149:15:@51011.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@51010.4]
  reg  regs_30; // @[SRAM.scala 145:20:@51017.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@51018.4]
  wire  _T_959; // @[SRAM.scala 148:25:@51019.4]
  wire  _T_960; // @[SRAM.scala 148:15:@51020.4]
  wire  _T_961; // @[SRAM.scala 149:15:@51022.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@51021.4]
  reg  regs_31; // @[SRAM.scala 145:20:@51028.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@51029.4]
  wire  _T_968; // @[SRAM.scala 148:25:@51030.4]
  wire  _T_969; // @[SRAM.scala 148:15:@51031.4]
  wire  _T_970; // @[SRAM.scala 149:15:@51033.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@51032.4]
  reg  regs_32; // @[SRAM.scala 145:20:@51039.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@51040.4]
  wire  _T_977; // @[SRAM.scala 148:25:@51041.4]
  wire  _T_978; // @[SRAM.scala 148:15:@51042.4]
  wire  _T_979; // @[SRAM.scala 149:15:@51044.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@51043.4]
  reg  regs_33; // @[SRAM.scala 145:20:@51050.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@51051.4]
  wire  _T_986; // @[SRAM.scala 148:25:@51052.4]
  wire  _T_987; // @[SRAM.scala 148:15:@51053.4]
  wire  _T_988; // @[SRAM.scala 149:15:@51055.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@51054.4]
  reg  regs_34; // @[SRAM.scala 145:20:@51061.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@51062.4]
  wire  _T_995; // @[SRAM.scala 148:25:@51063.4]
  wire  _T_996; // @[SRAM.scala 148:15:@51064.4]
  wire  _T_997; // @[SRAM.scala 149:15:@51066.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@51065.4]
  reg  regs_35; // @[SRAM.scala 145:20:@51072.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@51073.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@51074.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@51075.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@51077.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@51076.4]
  reg  regs_36; // @[SRAM.scala 145:20:@51083.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@51084.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@51085.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@51086.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@51088.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@51087.4]
  reg  regs_37; // @[SRAM.scala 145:20:@51094.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@51095.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@51096.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@51097.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@51099.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@51098.4]
  reg  regs_38; // @[SRAM.scala 145:20:@51105.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@51106.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@51107.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@51108.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@51110.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@51109.4]
  reg  regs_39; // @[SRAM.scala 145:20:@51116.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@51117.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@51118.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@51119.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@51121.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@51120.4]
  reg  regs_40; // @[SRAM.scala 145:20:@51127.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@51128.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@51129.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@51130.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@51132.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@51131.4]
  reg  regs_41; // @[SRAM.scala 145:20:@51138.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@51139.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@51140.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@51141.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@51143.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@51142.4]
  reg  regs_42; // @[SRAM.scala 145:20:@51149.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@51150.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@51151.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@51152.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@51154.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@51153.4]
  reg  regs_43; // @[SRAM.scala 145:20:@51160.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@51161.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@51162.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@51163.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@51165.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@51164.4]
  reg  regs_44; // @[SRAM.scala 145:20:@51171.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@51172.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@51173.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@51174.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@51176.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@51175.4]
  reg  regs_45; // @[SRAM.scala 145:20:@51182.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@51183.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@51184.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@51185.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@51187.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@51186.4]
  reg  regs_46; // @[SRAM.scala 145:20:@51193.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@51194.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@51195.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@51196.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@51198.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@51197.4]
  reg  regs_47; // @[SRAM.scala 145:20:@51204.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@51205.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@51206.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@51207.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@51209.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@51208.4]
  reg  regs_48; // @[SRAM.scala 145:20:@51215.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@51216.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@51217.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@51218.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@51220.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@51219.4]
  reg  regs_49; // @[SRAM.scala 145:20:@51226.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@51227.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@51228.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@51229.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@51231.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@51230.4]
  reg  regs_50; // @[SRAM.scala 145:20:@51237.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@51238.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@51239.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@51240.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@51242.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@51241.4]
  reg  regs_51; // @[SRAM.scala 145:20:@51248.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@51249.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@51250.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@51251.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@51253.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@51252.4]
  reg  regs_52; // @[SRAM.scala 145:20:@51259.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@51260.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@51261.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@51262.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@51264.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@51263.4]
  reg  regs_53; // @[SRAM.scala 145:20:@51270.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@51271.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@51272.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@51273.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@51275.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@51274.4]
  reg  regs_54; // @[SRAM.scala 145:20:@51281.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@51282.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@51283.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@51284.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@51286.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@51285.4]
  reg  regs_55; // @[SRAM.scala 145:20:@51292.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@51293.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@51294.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@51295.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@51297.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@51296.4]
  reg  regs_56; // @[SRAM.scala 145:20:@51303.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@51304.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@51305.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@51306.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@51308.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@51307.4]
  reg  regs_57; // @[SRAM.scala 145:20:@51314.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@51315.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@51316.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@51317.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@51319.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@51318.4]
  reg  regs_58; // @[SRAM.scala 145:20:@51325.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@51326.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@51327.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@51328.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@51330.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@51329.4]
  reg  regs_59; // @[SRAM.scala 145:20:@51336.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@51337.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@51338.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@51339.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@51341.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@51340.4]
  reg  regs_60; // @[SRAM.scala 145:20:@51347.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@51348.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@51349.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@51350.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@51352.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@51351.4]
  reg  regs_61; // @[SRAM.scala 145:20:@51358.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@51359.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@51360.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@51361.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@51363.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@51362.4]
  reg  regs_62; // @[SRAM.scala 145:20:@51369.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@51370.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@51371.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@51372.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@51374.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@51373.4]
  reg  regs_63; // @[SRAM.scala 145:20:@51380.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@51381.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@51382.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@51383.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@51385.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@51384.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@51454.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@51454.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@50688.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@50689.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@50690.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50692.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@50691.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@50699.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@50700.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@50701.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50703.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@50702.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@50710.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@50711.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@50712.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50714.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@50713.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@50721.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@50722.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@50723.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50725.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@50724.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@50732.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@50733.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@50734.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50736.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@50735.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@50743.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@50744.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@50745.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50747.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@50746.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@50754.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@50755.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@50756.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50758.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@50757.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@50765.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@50766.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@50767.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50769.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@50768.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@50776.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@50777.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@50778.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50780.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@50779.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@50787.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@50788.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@50789.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50791.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@50790.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@50798.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@50799.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@50800.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50802.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@50801.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@50809.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@50810.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@50811.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50813.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@50812.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@50820.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@50821.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@50822.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50824.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@50823.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@50831.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@50832.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@50833.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50835.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@50834.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@50842.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@50843.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@50844.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50846.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@50845.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@50853.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@50854.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@50855.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50857.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@50856.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@50864.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@50865.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@50866.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50868.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@50867.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@50875.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@50876.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@50877.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50879.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@50878.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@50886.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@50887.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@50888.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50890.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@50889.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@50897.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@50898.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@50899.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50901.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@50900.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@50908.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@50909.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@50910.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50912.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@50911.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@50919.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@50920.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@50921.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50923.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@50922.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@50930.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@50931.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@50932.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50934.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@50933.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@50941.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@50942.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@50943.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50945.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@50944.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@50952.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@50953.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@50954.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50956.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@50955.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@50963.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@50964.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@50965.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50967.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@50966.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@50974.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@50975.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@50976.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50978.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@50977.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@50985.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@50986.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@50987.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50989.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@50988.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@50996.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@50997.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@50998.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51000.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@50999.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@51007.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@51008.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@51009.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51011.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@51010.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@51018.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@51019.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@51020.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51022.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@51021.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@51029.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@51030.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@51031.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51033.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@51032.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@51040.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@51041.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@51042.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51044.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@51043.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@51051.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@51052.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@51053.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51055.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@51054.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@51062.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@51063.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@51064.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51066.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@51065.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@51073.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@51074.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@51075.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51077.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@51076.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@51084.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@51085.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@51086.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51088.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@51087.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@51095.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@51096.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@51097.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51099.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@51098.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@51106.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@51107.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@51108.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51110.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@51109.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@51117.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@51118.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@51119.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51121.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@51120.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@51128.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@51129.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@51130.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51132.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@51131.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@51139.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@51140.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@51141.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51143.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@51142.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@51150.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@51151.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@51152.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51154.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@51153.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@51161.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@51162.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@51163.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51165.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@51164.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@51172.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@51173.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@51174.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51176.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@51175.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@51183.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@51184.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@51185.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51187.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@51186.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@51194.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@51195.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@51196.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51198.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@51197.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@51205.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@51206.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@51207.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51209.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@51208.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@51216.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@51217.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@51218.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51220.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@51219.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@51227.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@51228.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@51229.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51231.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@51230.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@51238.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@51239.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@51240.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51242.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@51241.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@51249.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@51250.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@51251.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51253.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@51252.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@51260.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@51261.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@51262.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51264.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@51263.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@51271.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@51272.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@51273.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51275.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@51274.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@51282.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@51283.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@51284.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51286.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@51285.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@51293.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@51294.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@51295.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51297.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@51296.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@51304.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@51305.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@51306.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51308.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@51307.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@51315.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@51316.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@51317.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51319.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@51318.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@51326.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@51327.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@51328.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51330.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@51329.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@51337.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@51338.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@51339.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51341.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@51340.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@51348.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@51349.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@51350.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51352.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@51351.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@51359.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@51360.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@51361.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51363.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@51362.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@51370.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@51371.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@51372.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51374.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@51373.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@51381.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@51382.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@51383.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51385.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@51384.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@51454.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@51454.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@51454.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@51456.2]
  input   clock, // @[:@51457.4]
  input   reset, // @[:@51458.4]
  output  io_in_ready, // @[:@51459.4]
  input   io_in_valid, // @[:@51459.4]
  input   io_in_bits, // @[:@51459.4]
  input   io_out_ready, // @[:@51459.4]
  output  io_out_valid, // @[:@51459.4]
  output  io_out_bits, // @[:@51459.4]
  input   io_banks_0_wdata_valid, // @[:@51459.4]
  input   io_banks_0_wdata_bits, // @[:@51459.4]
  input   io_banks_1_wdata_valid, // @[:@51459.4]
  input   io_banks_1_wdata_bits, // @[:@51459.4]
  input   io_banks_2_wdata_valid, // @[:@51459.4]
  input   io_banks_2_wdata_bits, // @[:@51459.4]
  input   io_banks_3_wdata_valid, // @[:@51459.4]
  input   io_banks_3_wdata_bits, // @[:@51459.4]
  input   io_banks_4_wdata_valid, // @[:@51459.4]
  input   io_banks_4_wdata_bits, // @[:@51459.4]
  input   io_banks_5_wdata_valid, // @[:@51459.4]
  input   io_banks_5_wdata_bits, // @[:@51459.4]
  input   io_banks_6_wdata_valid, // @[:@51459.4]
  input   io_banks_6_wdata_bits, // @[:@51459.4]
  input   io_banks_7_wdata_valid, // @[:@51459.4]
  input   io_banks_7_wdata_bits, // @[:@51459.4]
  input   io_banks_8_wdata_valid, // @[:@51459.4]
  input   io_banks_8_wdata_bits, // @[:@51459.4]
  input   io_banks_9_wdata_valid, // @[:@51459.4]
  input   io_banks_9_wdata_bits, // @[:@51459.4]
  input   io_banks_10_wdata_valid, // @[:@51459.4]
  input   io_banks_10_wdata_bits, // @[:@51459.4]
  input   io_banks_11_wdata_valid, // @[:@51459.4]
  input   io_banks_11_wdata_bits, // @[:@51459.4]
  input   io_banks_12_wdata_valid, // @[:@51459.4]
  input   io_banks_12_wdata_bits, // @[:@51459.4]
  input   io_banks_13_wdata_valid, // @[:@51459.4]
  input   io_banks_13_wdata_bits, // @[:@51459.4]
  input   io_banks_14_wdata_valid, // @[:@51459.4]
  input   io_banks_14_wdata_bits, // @[:@51459.4]
  input   io_banks_15_wdata_valid, // @[:@51459.4]
  input   io_banks_15_wdata_bits, // @[:@51459.4]
  input   io_banks_16_wdata_valid, // @[:@51459.4]
  input   io_banks_16_wdata_bits, // @[:@51459.4]
  input   io_banks_17_wdata_valid, // @[:@51459.4]
  input   io_banks_17_wdata_bits, // @[:@51459.4]
  input   io_banks_18_wdata_valid, // @[:@51459.4]
  input   io_banks_18_wdata_bits, // @[:@51459.4]
  input   io_banks_19_wdata_valid, // @[:@51459.4]
  input   io_banks_19_wdata_bits, // @[:@51459.4]
  input   io_banks_20_wdata_valid, // @[:@51459.4]
  input   io_banks_20_wdata_bits, // @[:@51459.4]
  input   io_banks_21_wdata_valid, // @[:@51459.4]
  input   io_banks_21_wdata_bits, // @[:@51459.4]
  input   io_banks_22_wdata_valid, // @[:@51459.4]
  input   io_banks_22_wdata_bits, // @[:@51459.4]
  input   io_banks_23_wdata_valid, // @[:@51459.4]
  input   io_banks_23_wdata_bits, // @[:@51459.4]
  input   io_banks_24_wdata_valid, // @[:@51459.4]
  input   io_banks_24_wdata_bits, // @[:@51459.4]
  input   io_banks_25_wdata_valid, // @[:@51459.4]
  input   io_banks_25_wdata_bits, // @[:@51459.4]
  input   io_banks_26_wdata_valid, // @[:@51459.4]
  input   io_banks_26_wdata_bits, // @[:@51459.4]
  input   io_banks_27_wdata_valid, // @[:@51459.4]
  input   io_banks_27_wdata_bits, // @[:@51459.4]
  input   io_banks_28_wdata_valid, // @[:@51459.4]
  input   io_banks_28_wdata_bits, // @[:@51459.4]
  input   io_banks_29_wdata_valid, // @[:@51459.4]
  input   io_banks_29_wdata_bits, // @[:@51459.4]
  input   io_banks_30_wdata_valid, // @[:@51459.4]
  input   io_banks_30_wdata_bits, // @[:@51459.4]
  input   io_banks_31_wdata_valid, // @[:@51459.4]
  input   io_banks_31_wdata_bits, // @[:@51459.4]
  input   io_banks_32_wdata_valid, // @[:@51459.4]
  input   io_banks_32_wdata_bits, // @[:@51459.4]
  input   io_banks_33_wdata_valid, // @[:@51459.4]
  input   io_banks_33_wdata_bits, // @[:@51459.4]
  input   io_banks_34_wdata_valid, // @[:@51459.4]
  input   io_banks_34_wdata_bits, // @[:@51459.4]
  input   io_banks_35_wdata_valid, // @[:@51459.4]
  input   io_banks_35_wdata_bits, // @[:@51459.4]
  input   io_banks_36_wdata_valid, // @[:@51459.4]
  input   io_banks_36_wdata_bits, // @[:@51459.4]
  input   io_banks_37_wdata_valid, // @[:@51459.4]
  input   io_banks_37_wdata_bits, // @[:@51459.4]
  input   io_banks_38_wdata_valid, // @[:@51459.4]
  input   io_banks_38_wdata_bits, // @[:@51459.4]
  input   io_banks_39_wdata_valid, // @[:@51459.4]
  input   io_banks_39_wdata_bits, // @[:@51459.4]
  input   io_banks_40_wdata_valid, // @[:@51459.4]
  input   io_banks_40_wdata_bits, // @[:@51459.4]
  input   io_banks_41_wdata_valid, // @[:@51459.4]
  input   io_banks_41_wdata_bits, // @[:@51459.4]
  input   io_banks_42_wdata_valid, // @[:@51459.4]
  input   io_banks_42_wdata_bits, // @[:@51459.4]
  input   io_banks_43_wdata_valid, // @[:@51459.4]
  input   io_banks_43_wdata_bits, // @[:@51459.4]
  input   io_banks_44_wdata_valid, // @[:@51459.4]
  input   io_banks_44_wdata_bits, // @[:@51459.4]
  input   io_banks_45_wdata_valid, // @[:@51459.4]
  input   io_banks_45_wdata_bits, // @[:@51459.4]
  input   io_banks_46_wdata_valid, // @[:@51459.4]
  input   io_banks_46_wdata_bits, // @[:@51459.4]
  input   io_banks_47_wdata_valid, // @[:@51459.4]
  input   io_banks_47_wdata_bits, // @[:@51459.4]
  input   io_banks_48_wdata_valid, // @[:@51459.4]
  input   io_banks_48_wdata_bits, // @[:@51459.4]
  input   io_banks_49_wdata_valid, // @[:@51459.4]
  input   io_banks_49_wdata_bits, // @[:@51459.4]
  input   io_banks_50_wdata_valid, // @[:@51459.4]
  input   io_banks_50_wdata_bits, // @[:@51459.4]
  input   io_banks_51_wdata_valid, // @[:@51459.4]
  input   io_banks_51_wdata_bits, // @[:@51459.4]
  input   io_banks_52_wdata_valid, // @[:@51459.4]
  input   io_banks_52_wdata_bits, // @[:@51459.4]
  input   io_banks_53_wdata_valid, // @[:@51459.4]
  input   io_banks_53_wdata_bits, // @[:@51459.4]
  input   io_banks_54_wdata_valid, // @[:@51459.4]
  input   io_banks_54_wdata_bits, // @[:@51459.4]
  input   io_banks_55_wdata_valid, // @[:@51459.4]
  input   io_banks_55_wdata_bits, // @[:@51459.4]
  input   io_banks_56_wdata_valid, // @[:@51459.4]
  input   io_banks_56_wdata_bits, // @[:@51459.4]
  input   io_banks_57_wdata_valid, // @[:@51459.4]
  input   io_banks_57_wdata_bits, // @[:@51459.4]
  input   io_banks_58_wdata_valid, // @[:@51459.4]
  input   io_banks_58_wdata_bits, // @[:@51459.4]
  input   io_banks_59_wdata_valid, // @[:@51459.4]
  input   io_banks_59_wdata_bits, // @[:@51459.4]
  input   io_banks_60_wdata_valid, // @[:@51459.4]
  input   io_banks_60_wdata_bits, // @[:@51459.4]
  input   io_banks_61_wdata_valid, // @[:@51459.4]
  input   io_banks_61_wdata_bits, // @[:@51459.4]
  input   io_banks_62_wdata_valid, // @[:@51459.4]
  input   io_banks_62_wdata_bits, // @[:@51459.4]
  input   io_banks_63_wdata_valid, // @[:@51459.4]
  input   io_banks_63_wdata_bits // @[:@51459.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@51725.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@51725.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@51725.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@51725.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@51725.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@51735.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@51735.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@51735.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@51735.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@51735.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@51750.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@51750.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@51750.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@51750.4]
  wire  writeEn; // @[FIFO.scala 30:29:@51723.4]
  wire  readEn; // @[FIFO.scala 31:29:@51724.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@51745.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@51746.4]
  wire  _T_824; // @[FIFO.scala 45:27:@51747.4]
  wire  empty; // @[FIFO.scala 45:24:@51748.4]
  wire  full; // @[FIFO.scala 46:23:@51749.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@52916.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@52917.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@51725.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@51735.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@51750.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@51723.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@51724.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@51746.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@51747.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@51748.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@51749.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@52916.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@52917.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@52923.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@52921.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@51955.4]
  assign enqCounter_clock = clock; // @[:@51726.4]
  assign enqCounter_reset = reset; // @[:@51727.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@51733.4]
  assign deqCounter_clock = clock; // @[:@51736.4]
  assign deqCounter_reset = reset; // @[:@51737.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@51743.4]
  assign FFRAM_clock = clock; // @[:@51751.4]
  assign FFRAM_reset = reset; // @[:@51752.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@51951.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@51952.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@51953.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@51954.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@51957.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@51956.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@51960.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@51959.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@51963.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@51962.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@51966.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@51965.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@51969.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@51968.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@51972.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@51971.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@51975.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@51974.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@51978.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@51977.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@51981.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@51980.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@51984.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@51983.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@51987.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@51986.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@51990.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@51989.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@51993.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@51992.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@51996.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@51995.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@51999.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@51998.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@52002.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@52001.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@52005.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@52004.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@52008.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@52007.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@52011.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@52010.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@52014.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@52013.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@52017.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@52016.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@52020.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@52019.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@52023.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@52022.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@52026.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@52025.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@52029.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@52028.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@52032.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@52031.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@52035.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@52034.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@52038.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@52037.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@52041.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@52040.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@52044.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@52043.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@52047.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@52046.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@52050.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@52049.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@52053.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@52052.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@52056.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@52055.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@52059.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@52058.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@52062.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@52061.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@52065.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@52064.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@52068.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@52067.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@52071.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@52070.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@52074.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@52073.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@52077.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@52076.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@52080.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@52079.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@52083.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@52082.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@52086.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@52085.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@52089.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@52088.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@52092.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@52091.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@52095.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@52094.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@52098.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@52097.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@52101.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@52100.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@52104.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@52103.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@52107.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@52106.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@52110.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@52109.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@52113.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@52112.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@52116.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@52115.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@52119.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@52118.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@52122.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@52121.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@52125.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@52124.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@52128.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@52127.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@52131.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@52130.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@52134.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@52133.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@52137.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@52136.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@52140.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@52139.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@52143.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@52142.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@52146.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@52145.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@52925.2]
  input         clock, // @[:@52926.4]
  input         reset, // @[:@52927.4]
  input         io_dram_cmd_ready, // @[:@52928.4]
  output        io_dram_cmd_valid, // @[:@52928.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@52928.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@52928.4]
  input         io_dram_wdata_ready, // @[:@52928.4]
  output        io_dram_wdata_valid, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@52928.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@52928.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@52928.4]
  output        io_dram_wresp_ready, // @[:@52928.4]
  input         io_dram_wresp_valid, // @[:@52928.4]
  output        io_store_cmd_ready, // @[:@52928.4]
  input         io_store_cmd_valid, // @[:@52928.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@52928.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@52928.4]
  output        io_store_data_ready, // @[:@52928.4]
  input         io_store_data_valid, // @[:@52928.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@52928.4]
  input         io_store_data_bits_wstrb, // @[:@52928.4]
  input         io_store_wresp_ready, // @[:@52928.4]
  output        io_store_wresp_valid, // @[:@52928.4]
  output        io_store_wresp_bits // @[:@52928.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@53053.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@53053.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@53053.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@53053.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@53053.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@53053.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@53053.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@53053.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@53053.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@53053.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@53459.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@53459.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@53459.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@53459.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@53459.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@53459.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@53459.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@53459.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@53459.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@53700.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@53700.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@53456.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@53053.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@53459.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@53700.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@53456.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@53453.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@53454.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@53457.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@53489.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@53490.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@53491.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@53492.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@53493.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@53494.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@53495.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@53496.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@53497.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@53498.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@53499.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@53500.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@53501.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@53502.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@53503.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@53504.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@53505.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@53635.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@53636.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@53637.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@53638.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@53639.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@53640.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@53641.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@53642.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@53643.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@53644.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@53645.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@53646.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@53647.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@53648.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@53649.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@53650.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@53651.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@53652.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@53653.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@53654.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@53655.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@53656.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@53657.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@53658.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@53659.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@53660.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@53661.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@53662.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@53663.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@53664.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@53665.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@53666.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@53667.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@53668.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@53669.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@53670.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@53671.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@53672.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@53673.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@53674.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@53675.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@53676.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@53677.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@53678.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@53679.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@53680.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@53681.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@53682.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@53683.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@53684.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@53685.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@53686.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@53687.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@53688.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@53689.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@53690.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@53691.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@53692.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@53693.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@53694.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@53695.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@53696.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@53697.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@53698.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@53967.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@53451.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@53488.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@53968.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@53969.4]
  assign cmd_clock = clock; // @[:@53054.4]
  assign cmd_reset = reset; // @[:@53055.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@53448.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@53450.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@53449.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@53452.4]
  assign wdata_clock = clock; // @[:@53460.4]
  assign wdata_reset = reset; // @[:@53461.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@53485.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@53486.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@53487.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@53699.4]
  assign wresp_clock = clock; // @[:@53701.4]
  assign wresp_reset = reset; // @[:@53702.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@53965.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@53966.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@53970.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@54036.2]
  output        io_in_ready, // @[:@54039.4]
  input         io_in_valid, // @[:@54039.4]
  input  [63:0] io_in_bits_0_addr, // @[:@54039.4]
  input  [31:0] io_in_bits_0_size, // @[:@54039.4]
  input         io_in_bits_0_isWr, // @[:@54039.4]
  input  [31:0] io_in_bits_0_tag, // @[:@54039.4]
  input         io_out_ready, // @[:@54039.4]
  output        io_out_valid, // @[:@54039.4]
  output [63:0] io_out_bits_addr, // @[:@54039.4]
  output [31:0] io_out_bits_size, // @[:@54039.4]
  output        io_out_bits_isWr, // @[:@54039.4]
  output [31:0] io_out_bits_tag // @[:@54039.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@54041.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@54041.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@54050.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@54049.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@54055.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@54054.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@54052.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@54051.4]
endmodule
module MuxPipe_1( // @[:@54057.2]
  output        io_in_ready, // @[:@54060.4]
  input         io_in_valid, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@54060.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@54060.4]
  input         io_in_bits_0_wstrb_0, // @[:@54060.4]
  input         io_in_bits_0_wstrb_1, // @[:@54060.4]
  input         io_in_bits_0_wstrb_2, // @[:@54060.4]
  input         io_in_bits_0_wstrb_3, // @[:@54060.4]
  input         io_in_bits_0_wstrb_4, // @[:@54060.4]
  input         io_in_bits_0_wstrb_5, // @[:@54060.4]
  input         io_in_bits_0_wstrb_6, // @[:@54060.4]
  input         io_in_bits_0_wstrb_7, // @[:@54060.4]
  input         io_in_bits_0_wstrb_8, // @[:@54060.4]
  input         io_in_bits_0_wstrb_9, // @[:@54060.4]
  input         io_in_bits_0_wstrb_10, // @[:@54060.4]
  input         io_in_bits_0_wstrb_11, // @[:@54060.4]
  input         io_in_bits_0_wstrb_12, // @[:@54060.4]
  input         io_in_bits_0_wstrb_13, // @[:@54060.4]
  input         io_in_bits_0_wstrb_14, // @[:@54060.4]
  input         io_in_bits_0_wstrb_15, // @[:@54060.4]
  input         io_in_bits_0_wstrb_16, // @[:@54060.4]
  input         io_in_bits_0_wstrb_17, // @[:@54060.4]
  input         io_in_bits_0_wstrb_18, // @[:@54060.4]
  input         io_in_bits_0_wstrb_19, // @[:@54060.4]
  input         io_in_bits_0_wstrb_20, // @[:@54060.4]
  input         io_in_bits_0_wstrb_21, // @[:@54060.4]
  input         io_in_bits_0_wstrb_22, // @[:@54060.4]
  input         io_in_bits_0_wstrb_23, // @[:@54060.4]
  input         io_in_bits_0_wstrb_24, // @[:@54060.4]
  input         io_in_bits_0_wstrb_25, // @[:@54060.4]
  input         io_in_bits_0_wstrb_26, // @[:@54060.4]
  input         io_in_bits_0_wstrb_27, // @[:@54060.4]
  input         io_in_bits_0_wstrb_28, // @[:@54060.4]
  input         io_in_bits_0_wstrb_29, // @[:@54060.4]
  input         io_in_bits_0_wstrb_30, // @[:@54060.4]
  input         io_in_bits_0_wstrb_31, // @[:@54060.4]
  input         io_in_bits_0_wstrb_32, // @[:@54060.4]
  input         io_in_bits_0_wstrb_33, // @[:@54060.4]
  input         io_in_bits_0_wstrb_34, // @[:@54060.4]
  input         io_in_bits_0_wstrb_35, // @[:@54060.4]
  input         io_in_bits_0_wstrb_36, // @[:@54060.4]
  input         io_in_bits_0_wstrb_37, // @[:@54060.4]
  input         io_in_bits_0_wstrb_38, // @[:@54060.4]
  input         io_in_bits_0_wstrb_39, // @[:@54060.4]
  input         io_in_bits_0_wstrb_40, // @[:@54060.4]
  input         io_in_bits_0_wstrb_41, // @[:@54060.4]
  input         io_in_bits_0_wstrb_42, // @[:@54060.4]
  input         io_in_bits_0_wstrb_43, // @[:@54060.4]
  input         io_in_bits_0_wstrb_44, // @[:@54060.4]
  input         io_in_bits_0_wstrb_45, // @[:@54060.4]
  input         io_in_bits_0_wstrb_46, // @[:@54060.4]
  input         io_in_bits_0_wstrb_47, // @[:@54060.4]
  input         io_in_bits_0_wstrb_48, // @[:@54060.4]
  input         io_in_bits_0_wstrb_49, // @[:@54060.4]
  input         io_in_bits_0_wstrb_50, // @[:@54060.4]
  input         io_in_bits_0_wstrb_51, // @[:@54060.4]
  input         io_in_bits_0_wstrb_52, // @[:@54060.4]
  input         io_in_bits_0_wstrb_53, // @[:@54060.4]
  input         io_in_bits_0_wstrb_54, // @[:@54060.4]
  input         io_in_bits_0_wstrb_55, // @[:@54060.4]
  input         io_in_bits_0_wstrb_56, // @[:@54060.4]
  input         io_in_bits_0_wstrb_57, // @[:@54060.4]
  input         io_in_bits_0_wstrb_58, // @[:@54060.4]
  input         io_in_bits_0_wstrb_59, // @[:@54060.4]
  input         io_in_bits_0_wstrb_60, // @[:@54060.4]
  input         io_in_bits_0_wstrb_61, // @[:@54060.4]
  input         io_in_bits_0_wstrb_62, // @[:@54060.4]
  input         io_in_bits_0_wstrb_63, // @[:@54060.4]
  input         io_out_ready, // @[:@54060.4]
  output        io_out_valid, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_0, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_1, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_2, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_3, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_4, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_5, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_6, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_7, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_8, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_9, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_10, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_11, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_12, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_13, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_14, // @[:@54060.4]
  output [31:0] io_out_bits_wdata_15, // @[:@54060.4]
  output        io_out_bits_wstrb_0, // @[:@54060.4]
  output        io_out_bits_wstrb_1, // @[:@54060.4]
  output        io_out_bits_wstrb_2, // @[:@54060.4]
  output        io_out_bits_wstrb_3, // @[:@54060.4]
  output        io_out_bits_wstrb_4, // @[:@54060.4]
  output        io_out_bits_wstrb_5, // @[:@54060.4]
  output        io_out_bits_wstrb_6, // @[:@54060.4]
  output        io_out_bits_wstrb_7, // @[:@54060.4]
  output        io_out_bits_wstrb_8, // @[:@54060.4]
  output        io_out_bits_wstrb_9, // @[:@54060.4]
  output        io_out_bits_wstrb_10, // @[:@54060.4]
  output        io_out_bits_wstrb_11, // @[:@54060.4]
  output        io_out_bits_wstrb_12, // @[:@54060.4]
  output        io_out_bits_wstrb_13, // @[:@54060.4]
  output        io_out_bits_wstrb_14, // @[:@54060.4]
  output        io_out_bits_wstrb_15, // @[:@54060.4]
  output        io_out_bits_wstrb_16, // @[:@54060.4]
  output        io_out_bits_wstrb_17, // @[:@54060.4]
  output        io_out_bits_wstrb_18, // @[:@54060.4]
  output        io_out_bits_wstrb_19, // @[:@54060.4]
  output        io_out_bits_wstrb_20, // @[:@54060.4]
  output        io_out_bits_wstrb_21, // @[:@54060.4]
  output        io_out_bits_wstrb_22, // @[:@54060.4]
  output        io_out_bits_wstrb_23, // @[:@54060.4]
  output        io_out_bits_wstrb_24, // @[:@54060.4]
  output        io_out_bits_wstrb_25, // @[:@54060.4]
  output        io_out_bits_wstrb_26, // @[:@54060.4]
  output        io_out_bits_wstrb_27, // @[:@54060.4]
  output        io_out_bits_wstrb_28, // @[:@54060.4]
  output        io_out_bits_wstrb_29, // @[:@54060.4]
  output        io_out_bits_wstrb_30, // @[:@54060.4]
  output        io_out_bits_wstrb_31, // @[:@54060.4]
  output        io_out_bits_wstrb_32, // @[:@54060.4]
  output        io_out_bits_wstrb_33, // @[:@54060.4]
  output        io_out_bits_wstrb_34, // @[:@54060.4]
  output        io_out_bits_wstrb_35, // @[:@54060.4]
  output        io_out_bits_wstrb_36, // @[:@54060.4]
  output        io_out_bits_wstrb_37, // @[:@54060.4]
  output        io_out_bits_wstrb_38, // @[:@54060.4]
  output        io_out_bits_wstrb_39, // @[:@54060.4]
  output        io_out_bits_wstrb_40, // @[:@54060.4]
  output        io_out_bits_wstrb_41, // @[:@54060.4]
  output        io_out_bits_wstrb_42, // @[:@54060.4]
  output        io_out_bits_wstrb_43, // @[:@54060.4]
  output        io_out_bits_wstrb_44, // @[:@54060.4]
  output        io_out_bits_wstrb_45, // @[:@54060.4]
  output        io_out_bits_wstrb_46, // @[:@54060.4]
  output        io_out_bits_wstrb_47, // @[:@54060.4]
  output        io_out_bits_wstrb_48, // @[:@54060.4]
  output        io_out_bits_wstrb_49, // @[:@54060.4]
  output        io_out_bits_wstrb_50, // @[:@54060.4]
  output        io_out_bits_wstrb_51, // @[:@54060.4]
  output        io_out_bits_wstrb_52, // @[:@54060.4]
  output        io_out_bits_wstrb_53, // @[:@54060.4]
  output        io_out_bits_wstrb_54, // @[:@54060.4]
  output        io_out_bits_wstrb_55, // @[:@54060.4]
  output        io_out_bits_wstrb_56, // @[:@54060.4]
  output        io_out_bits_wstrb_57, // @[:@54060.4]
  output        io_out_bits_wstrb_58, // @[:@54060.4]
  output        io_out_bits_wstrb_59, // @[:@54060.4]
  output        io_out_bits_wstrb_60, // @[:@54060.4]
  output        io_out_bits_wstrb_61, // @[:@54060.4]
  output        io_out_bits_wstrb_62, // @[:@54060.4]
  output        io_out_bits_wstrb_63 // @[:@54060.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@54062.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@54062.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@54147.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@54146.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@54213.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@54214.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@54215.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@54216.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@54217.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@54218.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@54219.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@54220.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@54221.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@54222.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@54223.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@54224.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@54225.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@54226.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@54227.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@54228.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@54149.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@54150.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@54151.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@54152.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@54153.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@54154.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@54155.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@54156.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@54157.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@54158.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@54159.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@54160.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@54161.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@54162.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@54163.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@54164.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@54165.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@54166.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@54167.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@54168.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@54169.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@54170.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@54171.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@54172.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@54173.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@54174.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@54175.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@54176.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@54177.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@54178.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@54179.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@54180.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@54181.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@54182.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@54183.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@54184.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@54185.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@54186.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@54187.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@54188.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@54189.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@54190.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@54191.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@54192.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@54193.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@54194.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@54195.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@54196.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@54197.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@54198.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@54199.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@54200.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@54201.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@54202.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@54203.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@54204.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@54205.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@54206.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@54207.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@54208.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@54209.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@54210.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@54211.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@54212.4]
endmodule
module ElementCounter( // @[:@54230.2]
  input         clock, // @[:@54231.4]
  input         reset, // @[:@54232.4]
  input         io_reset, // @[:@54233.4]
  input         io_enable, // @[:@54233.4]
  output [31:0] io_out // @[:@54233.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@54235.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@54236.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@54237.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@54242.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@54238.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@54236.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@54237.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@54242.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@54238.4]
  assign io_out = count; // @[Counter.scala 47:10:@54245.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@54247.2]
  input         clock, // @[:@54248.4]
  input         reset, // @[:@54249.4]
  output        io_app_0_cmd_ready, // @[:@54250.4]
  input         io_app_0_cmd_valid, // @[:@54250.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@54250.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@54250.4]
  input         io_app_0_cmd_bits_isWr, // @[:@54250.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@54250.4]
  output        io_app_0_wdata_ready, // @[:@54250.4]
  input         io_app_0_wdata_valid, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@54250.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@54250.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@54250.4]
  input         io_app_0_rresp_ready, // @[:@54250.4]
  input         io_app_0_wresp_ready, // @[:@54250.4]
  output        io_app_0_wresp_valid, // @[:@54250.4]
  input         io_dram_cmd_ready, // @[:@54250.4]
  output        io_dram_cmd_valid, // @[:@54250.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@54250.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@54250.4]
  output        io_dram_cmd_bits_isWr, // @[:@54250.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@54250.4]
  input         io_dram_wdata_ready, // @[:@54250.4]
  output        io_dram_wdata_valid, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@54250.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@54250.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@54250.4]
  output        io_dram_rresp_ready, // @[:@54250.4]
  output        io_dram_wresp_ready, // @[:@54250.4]
  input         io_dram_wresp_valid, // @[:@54250.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@54250.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@54479.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@54479.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@54479.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@54479.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@54479.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@54486.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@54486.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@54486.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@54486.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@54486.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@54496.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@54496.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@54496.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@54496.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@54496.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@54496.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@54496.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@54496.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@54496.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@54496.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@54496.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@54496.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@54519.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@54519.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@54522.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@54522.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@54522.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@54522.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@54522.4]
  wire  _T_346; // @[package.scala 96:25:@54491.4 package.scala 96:25:@54492.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@54493.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@54495.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@54511.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@54513.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@54516.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@54525.4]
  wire [31:0] _T_365; // @[:@54529.4 :@54530.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@54531.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@54537.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@54540.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@54541.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@54728.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@54735.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@54740.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@54744.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@54745.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@54769.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@54479.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@54486.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@54496.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@54519.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@54522.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@54491.4 package.scala 96:25:@54492.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@54493.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@54495.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@54511.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@54513.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@54516.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@54525.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@54529.4 :@54530.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@54531.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@54537.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@54540.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@54541.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@54728.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@54735.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@54740.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@54744.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@54745.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@54769.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@54742.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@54748.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@54771.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@54631.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@54630.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@54629.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@54627.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@54626.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@54714.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@54698.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@54699.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@54700.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@54701.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@54702.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@54703.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@54704.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@54705.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@54706.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@54707.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@54708.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@54709.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@54710.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@54711.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@54712.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@54713.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@54634.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@54635.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@54636.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@54637.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@54638.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@54639.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@54640.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@54641.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@54642.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@54643.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@54644.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@54645.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@54646.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@54647.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@54648.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@54649.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@54650.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@54651.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@54652.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@54653.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@54654.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@54655.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@54656.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@54657.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@54658.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@54659.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@54660.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@54661.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@54662.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@54663.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@54664.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@54665.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@54666.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@54667.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@54668.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@54669.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@54670.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@54671.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@54672.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@54673.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@54674.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@54675.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@54676.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@54677.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@54678.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@54679.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@54680.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@54681.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@54682.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@54683.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@54684.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@54685.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@54686.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@54687.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@54688.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@54689.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@54690.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@54691.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@54692.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@54693.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@54694.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@54695.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@54696.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@54697.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@54775.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@54778.4]
  assign RetimeWrapper_clock = clock; // @[:@54480.4]
  assign RetimeWrapper_reset = reset; // @[:@54481.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@54483.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@54482.4]
  assign RetimeWrapper_1_clock = clock; // @[:@54487.4]
  assign RetimeWrapper_1_reset = reset; // @[:@54488.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@54490.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@54489.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@54499.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@54505.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@54504.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@54502.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@54501.4 FringeBundles.scala 115:32:@54518.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@54632.4 StreamArbiter.scala 57:23:@54738.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@54543.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@54610.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@54611.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@54612.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@54613.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@54614.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@54615.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@54616.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@54617.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@54618.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@54619.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@54620.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@54621.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@54622.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@54623.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@54624.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@54625.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@54546.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@54547.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@54548.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@54549.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@54550.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@54551.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@54552.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@54553.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@54554.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@54555.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@54556.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@54557.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@54558.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@54559.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@54560.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@54561.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@54562.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@54563.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@54564.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@54565.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@54566.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@54567.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@54568.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@54569.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@54570.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@54571.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@54572.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@54573.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@54574.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@54575.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@54576.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@54577.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@54578.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@54579.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@54580.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@54581.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@54582.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@54583.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@54584.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@54585.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@54586.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@54587.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@54588.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@54589.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@54590.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@54591.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@54592.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@54593.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@54594.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@54595.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@54596.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@54597.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@54598.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@54599.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@54600.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@54601.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@54602.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@54603.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@54604.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@54605.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@54606.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@54607.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@54608.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@54609.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@54715.4 StreamArbiter.scala 58:25:@54739.4]
  assign elementCtr_clock = clock; // @[:@54523.4]
  assign elementCtr_reset = reset; // @[:@54524.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@54527.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@54526.4]
endmodule
module Counter_72( // @[:@54780.2]
  input         clock, // @[:@54781.4]
  input         reset, // @[:@54782.4]
  input         io_reset, // @[:@54783.4]
  input         io_enable, // @[:@54783.4]
  input  [31:0] io_stride, // @[:@54783.4]
  output [31:0] io_out, // @[:@54783.4]
  output [31:0] io_next // @[:@54783.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@54785.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@54786.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@54787.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@54792.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@54788.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@54786.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@54787.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@54792.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@54788.4]
  assign io_out = count; // @[Counter.scala 25:10:@54795.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@54796.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@54798.2]
  input         clock, // @[:@54799.4]
  input         reset, // @[:@54800.4]
  output        io_in_cmd_ready, // @[:@54801.4]
  input         io_in_cmd_valid, // @[:@54801.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@54801.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@54801.4]
  input         io_in_cmd_bits_isWr, // @[:@54801.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@54801.4]
  output        io_in_wdata_ready, // @[:@54801.4]
  input         io_in_wdata_valid, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@54801.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@54801.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@54801.4]
  input         io_in_rresp_ready, // @[:@54801.4]
  input         io_in_wresp_ready, // @[:@54801.4]
  output        io_in_wresp_valid, // @[:@54801.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@54801.4]
  input         io_out_cmd_ready, // @[:@54801.4]
  output        io_out_cmd_valid, // @[:@54801.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@54801.4]
  output [31:0] io_out_cmd_bits_size, // @[:@54801.4]
  output        io_out_cmd_bits_isWr, // @[:@54801.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@54801.4]
  input         io_out_wdata_ready, // @[:@54801.4]
  output        io_out_wdata_valid, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@54801.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@54801.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@54801.4]
  output        io_out_rresp_ready, // @[:@54801.4]
  output        io_out_wresp_ready, // @[:@54801.4]
  input         io_out_wresp_valid, // @[:@54801.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@54801.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@54915.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@54915.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@54915.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@54915.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@54915.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@54915.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@54915.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@54918.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@54919.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@54920.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@54921.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@54924.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@54924.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@54925.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@54925.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@54926.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@54929.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@54936.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@54940.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@54943.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@54946.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@54957.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@54915.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@54918.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@54919.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@54920.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@54921.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@54924.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@54924.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@54925.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@54925.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@54926.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@54929.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@54936.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@54940.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@54943.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@54946.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@54957.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@54914.4 AXIProtocol.scala 38:19:@54948.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@54907.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@54804.4 AXIProtocol.scala 46:21:@54962.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@54803.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@54913.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@54912.4 AXIProtocol.scala 29:24:@54931.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@54911.4 AXIProtocol.scala 25:24:@54923.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@54909.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@54908.4 FringeBundles.scala 115:32:@54945.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@54906.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@54890.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@54891.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@54892.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@54893.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@54894.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@54895.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@54896.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@54897.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@54898.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@54899.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@54900.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@54901.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@54902.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@54903.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@54904.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@54905.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@54826.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@54827.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@54828.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@54829.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@54830.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@54831.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@54832.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@54833.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@54834.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@54835.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@54836.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@54837.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@54838.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@54839.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@54840.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@54841.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@54842.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@54843.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@54844.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@54845.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@54846.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@54847.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@54848.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@54849.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@54850.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@54851.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@54852.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@54853.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@54854.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@54855.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@54856.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@54857.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@54858.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@54859.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@54860.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@54861.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@54862.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@54863.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@54864.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@54865.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@54866.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@54867.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@54868.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@54869.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@54870.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@54871.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@54872.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@54873.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@54874.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@54875.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@54876.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@54877.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@54878.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@54879.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@54880.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@54881.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@54882.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@54883.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@54884.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@54885.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@54886.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@54887.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@54888.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@54889.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@54824.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@54805.4 AXIProtocol.scala 47:22:@54964.4]
  assign cmdSizeCounter_clock = clock; // @[:@54916.4]
  assign cmdSizeCounter_reset = reset; // @[:@54917.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@54949.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@54950.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@54951.4]
endmodule
module AXICmdIssue( // @[:@54984.2]
  input         clock, // @[:@54985.4]
  input         reset, // @[:@54986.4]
  output        io_in_cmd_ready, // @[:@54987.4]
  input         io_in_cmd_valid, // @[:@54987.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@54987.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@54987.4]
  input         io_in_cmd_bits_isWr, // @[:@54987.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@54987.4]
  output        io_in_wdata_ready, // @[:@54987.4]
  input         io_in_wdata_valid, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@54987.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@54987.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@54987.4]
  input         io_in_rresp_ready, // @[:@54987.4]
  input         io_in_wresp_ready, // @[:@54987.4]
  output        io_in_wresp_valid, // @[:@54987.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@54987.4]
  input         io_out_cmd_ready, // @[:@54987.4]
  output        io_out_cmd_valid, // @[:@54987.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@54987.4]
  output [31:0] io_out_cmd_bits_size, // @[:@54987.4]
  output        io_out_cmd_bits_isWr, // @[:@54987.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@54987.4]
  input         io_out_wdata_ready, // @[:@54987.4]
  output        io_out_wdata_valid, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@54987.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@54987.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@54987.4]
  output        io_out_wdata_bits_wlast, // @[:@54987.4]
  output        io_out_rresp_ready, // @[:@54987.4]
  output        io_out_wresp_ready, // @[:@54987.4]
  input         io_out_wresp_valid, // @[:@54987.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@54987.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@55101.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@55101.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@55101.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@55101.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@55101.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@55101.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@55101.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@55104.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@55105.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@55106.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@55107.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@55108.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@55114.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@55115.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@55110.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@55124.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@55125.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@55101.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@55105.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@55106.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@55107.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@55108.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@55114.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@55115.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@55110.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@55124.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@55125.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@55100.4 AXIProtocol.scala 81:19:@55122.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@55093.4 AXIProtocol.scala 82:21:@55123.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@54990.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@54989.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@55099.4 AXIProtocol.scala 84:20:@55127.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@55098.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@55097.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@55095.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@55094.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@55092.4 AXIProtocol.scala 86:22:@55129.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@55076.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@55077.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@55078.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@55079.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@55080.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@55081.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@55082.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@55083.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@55084.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@55085.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@55086.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@55087.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@55088.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@55089.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@55090.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@55091.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@55012.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@55013.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@55014.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@55015.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@55016.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@55017.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@55018.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@55019.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@55020.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@55021.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@55022.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@55023.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@55024.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@55025.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@55026.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@55027.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@55028.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@55029.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@55030.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@55031.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@55032.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@55033.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@55034.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@55035.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@55036.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@55037.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@55038.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@55039.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@55040.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@55041.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@55042.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@55043.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@55044.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@55045.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@55046.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@55047.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@55048.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@55049.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@55050.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@55051.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@55052.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@55053.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@55054.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@55055.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@55056.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@55057.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@55058.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@55059.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@55060.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@55061.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@55062.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@55063.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@55064.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@55065.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@55066.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@55067.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@55068.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@55069.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@55070.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@55071.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@55072.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@55073.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@55074.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@55075.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@55011.4 AXIProtocol.scala 87:27:@55130.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@55010.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@54991.4]
  assign wdataCounter_clock = clock; // @[:@55102.4]
  assign wdataCounter_reset = reset; // @[:@55103.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@55118.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@55119.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@55120.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@55132.2]
  input         clock, // @[:@55133.4]
  input         reset, // @[:@55134.4]
  input         io_enable, // @[:@55135.4]
  output        io_app_stores_0_cmd_ready, // @[:@55135.4]
  input         io_app_stores_0_cmd_valid, // @[:@55135.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@55135.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@55135.4]
  output        io_app_stores_0_data_ready, // @[:@55135.4]
  input         io_app_stores_0_data_valid, // @[:@55135.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@55135.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@55135.4]
  input         io_app_stores_0_wresp_ready, // @[:@55135.4]
  output        io_app_stores_0_wresp_valid, // @[:@55135.4]
  output        io_app_stores_0_wresp_bits, // @[:@55135.4]
  input         io_dram_cmd_ready, // @[:@55135.4]
  output        io_dram_cmd_valid, // @[:@55135.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@55135.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@55135.4]
  output        io_dram_cmd_bits_isWr, // @[:@55135.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@55135.4]
  input         io_dram_wdata_ready, // @[:@55135.4]
  output        io_dram_wdata_valid, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@55135.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@55135.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@55135.4]
  output        io_dram_wdata_bits_wlast, // @[:@55135.4]
  output        io_dram_rresp_ready, // @[:@55135.4]
  output        io_dram_wresp_ready, // @[:@55135.4]
  input         io_dram_wresp_valid, // @[:@55135.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@55135.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@56021.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@56035.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@56263.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@56378.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@56378.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@56021.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@56035.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@56263.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@56378.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@56034.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@56030.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@56025.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@56024.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@56603.4 DRAMArbiter.scala 100:23:@56606.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@56602.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@56601.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@56599.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@56598.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@56596.4 DRAMArbiter.scala 101:25:@56608.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@56580.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@56581.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@56582.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@56583.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@56584.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@56585.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@56586.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@56587.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@56588.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@56589.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@56590.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@56591.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@56592.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@56593.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@56594.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@56595.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@56516.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@56517.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@56518.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@56519.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@56520.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@56521.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@56522.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@56523.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@56524.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@56525.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@56526.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@56527.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@56528.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@56529.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@56530.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@56531.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@56532.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@56533.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@56534.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@56535.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@56536.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@56537.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@56538.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@56539.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@56540.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@56541.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@56542.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@56543.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@56544.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@56545.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@56546.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@56547.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@56548.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@56549.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@56550.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@56551.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@56552.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@56553.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@56554.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@56555.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@56556.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@56557.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@56558.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@56559.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@56560.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@56561.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@56562.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@56563.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@56564.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@56565.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@56566.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@56567.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@56568.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@56569.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@56570.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@56571.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@56572.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@56573.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@56574.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@56575.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@56576.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@56577.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@56578.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@56579.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@56515.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@56514.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@56495.4]
  assign StreamControllerStore_clock = clock; // @[:@56022.4]
  assign StreamControllerStore_reset = reset; // @[:@56023.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@56150.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@56143.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@56040.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@56033.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@56032.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@56031.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@56029.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@56028.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@56027.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@56026.4]
  assign StreamArbiter_clock = clock; // @[:@56036.4]
  assign StreamArbiter_reset = reset; // @[:@56037.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@56261.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@56260.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@56259.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@56257.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@56256.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@56254.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@56238.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@56239.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@56240.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@56241.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@56242.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@56243.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@56244.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@56245.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@56246.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@56247.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@56248.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@56249.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@56250.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@56251.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@56252.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@56253.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@56174.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@56175.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@56176.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@56177.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@56178.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@56179.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@56180.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@56181.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@56182.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@56183.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@56184.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@56185.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@56186.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@56187.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@56188.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@56189.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@56190.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@56191.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@56192.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@56193.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@56194.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@56195.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@56196.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@56197.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@56198.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@56199.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@56200.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@56201.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@56202.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@56203.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@56204.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@56205.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@56206.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@56207.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@56208.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@56209.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@56210.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@56211.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@56212.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@56213.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@56214.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@56215.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@56216.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@56217.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@56218.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@56219.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@56220.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@56221.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@56222.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@56223.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@56224.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@56225.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@56226.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@56227.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@56228.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@56229.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@56230.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@56231.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@56232.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@56233.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@56234.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@56235.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@56236.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@56237.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@56172.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@56153.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@56377.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@56370.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@56267.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@56266.4]
  assign AXICmdSplit_clock = clock; // @[:@56264.4]
  assign AXICmdSplit_reset = reset; // @[:@56265.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@56376.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@56375.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@56374.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@56372.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@56371.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@56369.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@56353.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@56354.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@56355.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@56356.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@56357.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@56358.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@56359.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@56360.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@56361.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@56362.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@56363.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@56364.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@56365.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@56366.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@56367.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@56368.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@56289.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@56290.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@56291.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@56292.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@56293.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@56294.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@56295.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@56296.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@56297.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@56298.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@56299.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@56300.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@56301.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@56302.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@56303.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@56304.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@56305.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@56306.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@56307.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@56308.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@56309.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@56310.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@56311.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@56312.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@56313.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@56314.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@56315.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@56316.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@56317.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@56318.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@56319.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@56320.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@56321.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@56322.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@56323.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@56324.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@56325.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@56326.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@56327.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@56328.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@56329.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@56330.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@56331.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@56332.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@56333.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@56334.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@56335.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@56336.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@56337.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@56338.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@56339.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@56340.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@56341.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@56342.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@56343.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@56344.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@56345.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@56346.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@56347.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@56348.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@56349.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@56350.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@56351.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@56352.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@56287.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@56268.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@56492.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@56485.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@56382.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@56381.4]
  assign AXICmdIssue_clock = clock; // @[:@56379.4]
  assign AXICmdIssue_reset = reset; // @[:@56380.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@56491.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@56490.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@56489.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@56487.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@56486.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@56484.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@56468.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@56469.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@56470.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@56471.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@56472.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@56473.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@56474.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@56475.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@56476.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@56477.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@56478.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@56479.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@56480.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@56481.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@56482.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@56483.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@56404.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@56405.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@56406.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@56407.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@56408.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@56409.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@56410.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@56411.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@56412.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@56413.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@56414.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@56415.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@56416.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@56417.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@56418.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@56419.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@56420.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@56421.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@56422.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@56423.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@56424.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@56425.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@56426.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@56427.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@56428.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@56429.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@56430.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@56431.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@56432.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@56433.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@56434.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@56435.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@56436.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@56437.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@56438.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@56439.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@56440.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@56441.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@56442.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@56443.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@56444.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@56445.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@56446.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@56447.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@56448.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@56449.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@56450.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@56451.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@56452.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@56453.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@56454.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@56455.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@56456.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@56457.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@56458.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@56459.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@56460.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@56461.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@56462.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@56463.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@56464.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@56465.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@56466.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@56467.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@56402.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@56383.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@56604.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@56597.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@56494.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@56493.4]
endmodule
module DRAMArbiter_1( // @[:@70833.2]
  input         clock, // @[:@70834.4]
  input         reset, // @[:@70835.4]
  input         io_enable, // @[:@70836.4]
  input         io_dram_cmd_ready, // @[:@70836.4]
  output        io_dram_cmd_valid, // @[:@70836.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@70836.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@70836.4]
  output        io_dram_cmd_bits_isWr, // @[:@70836.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@70836.4]
  input         io_dram_wdata_ready, // @[:@70836.4]
  output        io_dram_wdata_valid, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@70836.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@70836.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@70836.4]
  output        io_dram_wdata_bits_wlast, // @[:@70836.4]
  output        io_dram_rresp_ready, // @[:@70836.4]
  output        io_dram_wresp_ready, // @[:@70836.4]
  input         io_dram_wresp_valid, // @[:@70836.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@70836.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@71722.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@71736.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@71964.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@72079.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@72079.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@71722.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@71736.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@71964.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@72079.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@72304.4 DRAMArbiter.scala 100:23:@72307.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@72303.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@72302.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@72300.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@72299.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@72297.4 DRAMArbiter.scala 101:25:@72309.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@72281.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@72282.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@72283.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@72284.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@72285.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@72286.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@72287.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@72288.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@72289.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@72290.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@72291.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@72292.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@72293.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@72294.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@72295.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@72296.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@72217.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@72218.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@72219.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@72220.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@72221.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@72222.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@72223.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@72224.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@72225.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@72226.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@72227.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@72228.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@72229.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@72230.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@72231.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@72232.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@72233.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@72234.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@72235.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@72236.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@72237.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@72238.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@72239.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@72240.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@72241.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@72242.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@72243.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@72244.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@72245.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@72246.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@72247.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@72248.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@72249.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@72250.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@72251.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@72252.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@72253.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@72254.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@72255.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@72256.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@72257.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@72258.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@72259.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@72260.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@72261.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@72262.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@72263.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@72264.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@72265.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@72266.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@72267.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@72268.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@72269.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@72270.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@72271.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@72272.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@72273.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@72274.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@72275.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@72276.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@72277.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@72278.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@72279.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@72280.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@72216.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@72215.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@72196.4]
  assign StreamControllerStore_clock = clock; // @[:@71723.4]
  assign StreamControllerStore_reset = reset; // @[:@71724.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@71851.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@71844.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@71741.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@71734.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@71733.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@71732.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@71730.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@71729.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@71728.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@71727.4]
  assign StreamArbiter_clock = clock; // @[:@71737.4]
  assign StreamArbiter_reset = reset; // @[:@71738.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@71962.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@71961.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@71960.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@71958.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@71957.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@71955.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@71939.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@71940.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@71941.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@71942.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@71943.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@71944.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@71945.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@71946.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@71947.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@71948.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@71949.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@71950.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@71951.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@71952.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@71953.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@71954.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@71875.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@71876.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@71877.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@71878.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@71879.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@71880.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@71881.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@71882.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@71883.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@71884.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@71885.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@71886.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@71887.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@71888.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@71889.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@71890.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@71891.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@71892.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@71893.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@71894.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@71895.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@71896.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@71897.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@71898.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@71899.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@71900.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@71901.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@71902.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@71903.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@71904.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@71905.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@71906.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@71907.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@71908.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@71909.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@71910.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@71911.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@71912.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@71913.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@71914.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@71915.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@71916.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@71917.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@71918.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@71919.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@71920.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@71921.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@71922.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@71923.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@71924.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@71925.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@71926.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@71927.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@71928.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@71929.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@71930.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@71931.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@71932.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@71933.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@71934.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@71935.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@71936.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@71937.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@71938.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@71873.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@71854.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@72078.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@72071.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@71968.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@71967.4]
  assign AXICmdSplit_clock = clock; // @[:@71965.4]
  assign AXICmdSplit_reset = reset; // @[:@71966.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@72077.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@72076.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@72075.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@72073.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@72072.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@72070.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@72054.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@72055.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@72056.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@72057.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@72058.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@72059.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@72060.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@72061.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@72062.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@72063.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@72064.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@72065.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@72066.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@72067.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@72068.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@72069.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@71990.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@71991.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@71992.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@71993.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@71994.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@71995.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@71996.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@71997.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@71998.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@71999.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@72000.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@72001.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@72002.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@72003.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@72004.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@72005.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@72006.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@72007.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@72008.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@72009.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@72010.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@72011.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@72012.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@72013.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@72014.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@72015.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@72016.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@72017.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@72018.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@72019.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@72020.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@72021.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@72022.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@72023.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@72024.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@72025.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@72026.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@72027.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@72028.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@72029.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@72030.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@72031.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@72032.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@72033.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@72034.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@72035.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@72036.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@72037.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@72038.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@72039.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@72040.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@72041.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@72042.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@72043.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@72044.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@72045.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@72046.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@72047.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@72048.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@72049.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@72050.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@72051.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@72052.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@72053.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@71988.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@71969.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@72193.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@72186.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@72083.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@72082.4]
  assign AXICmdIssue_clock = clock; // @[:@72080.4]
  assign AXICmdIssue_reset = reset; // @[:@72081.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@72192.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@72191.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@72190.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@72188.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@72187.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@72185.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@72169.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@72170.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@72171.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@72172.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@72173.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@72174.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@72175.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@72176.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@72177.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@72178.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@72179.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@72180.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@72181.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@72182.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@72183.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@72184.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@72105.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@72106.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@72107.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@72108.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@72109.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@72110.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@72111.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@72112.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@72113.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@72114.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@72115.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@72116.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@72117.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@72118.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@72119.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@72120.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@72121.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@72122.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@72123.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@72124.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@72125.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@72126.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@72127.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@72128.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@72129.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@72130.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@72131.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@72132.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@72133.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@72134.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@72135.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@72136.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@72137.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@72138.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@72139.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@72140.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@72141.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@72142.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@72143.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@72144.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@72145.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@72146.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@72147.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@72148.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@72149.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@72150.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@72151.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@72152.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@72153.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@72154.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@72155.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@72156.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@72157.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@72158.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@72159.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@72160.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@72161.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@72162.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@72163.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@72164.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@72165.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@72166.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@72167.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@72168.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@72103.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@72084.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@72305.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@72298.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@72195.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@72194.4]
endmodule
module DRAMHeap( // @[:@102941.2]
  input         io_accel_0_req_valid, // @[:@102944.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@102944.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@102944.4]
  output        io_accel_0_resp_valid, // @[:@102944.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@102944.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@102944.4]
  output        io_host_0_req_valid, // @[:@102944.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@102944.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@102944.4]
  input         io_host_0_resp_valid, // @[:@102944.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@102944.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@102944.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@102951.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@102953.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@102952.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@102948.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@102947.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@102946.4]
endmodule
module RetimeWrapper_420( // @[:@102967.2]
  input         clock, // @[:@102968.4]
  input         reset, // @[:@102969.4]
  input         io_flow, // @[:@102970.4]
  input  [63:0] io_in, // @[:@102970.4]
  output [63:0] io_out // @[:@102970.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@102972.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@102972.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@102972.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@102972.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@102972.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@102972.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@102972.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@102985.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@102984.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@102983.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@102982.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@102981.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@102979.4]
endmodule
module FringeFF( // @[:@102987.2]
  input         clock, // @[:@102988.4]
  input         reset, // @[:@102989.4]
  input  [63:0] io_in, // @[:@102990.4]
  input         io_reset, // @[:@102990.4]
  output [63:0] io_out, // @[:@102990.4]
  input         io_enable // @[:@102990.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@102993.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@102993.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@102993.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@102993.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@102993.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@102998.4 package.scala 96:25:@102999.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@103004.6]
  RetimeWrapper_420 RetimeWrapper ( // @[package.scala 93:22:@102993.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@102998.4 package.scala 96:25:@102999.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@103004.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@103010.4]
  assign RetimeWrapper_clock = clock; // @[:@102994.4]
  assign RetimeWrapper_reset = reset; // @[:@102995.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@102997.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@102996.4]
endmodule
module MuxN( // @[:@131626.2]
  input  [63:0] io_ins_0, // @[:@131629.4]
  input  [63:0] io_ins_1, // @[:@131629.4]
  input  [63:0] io_ins_2, // @[:@131629.4]
  input  [63:0] io_ins_3, // @[:@131629.4]
  input  [63:0] io_ins_4, // @[:@131629.4]
  input  [63:0] io_ins_5, // @[:@131629.4]
  input  [63:0] io_ins_6, // @[:@131629.4]
  input  [63:0] io_ins_7, // @[:@131629.4]
  input  [63:0] io_ins_8, // @[:@131629.4]
  input  [63:0] io_ins_9, // @[:@131629.4]
  input  [63:0] io_ins_10, // @[:@131629.4]
  input  [63:0] io_ins_11, // @[:@131629.4]
  input  [63:0] io_ins_12, // @[:@131629.4]
  input  [63:0] io_ins_13, // @[:@131629.4]
  input  [63:0] io_ins_14, // @[:@131629.4]
  input  [63:0] io_ins_15, // @[:@131629.4]
  input  [63:0] io_ins_16, // @[:@131629.4]
  input  [63:0] io_ins_17, // @[:@131629.4]
  input  [63:0] io_ins_18, // @[:@131629.4]
  input  [63:0] io_ins_19, // @[:@131629.4]
  input  [63:0] io_ins_20, // @[:@131629.4]
  input  [63:0] io_ins_21, // @[:@131629.4]
  input  [63:0] io_ins_22, // @[:@131629.4]
  input  [63:0] io_ins_23, // @[:@131629.4]
  input  [63:0] io_ins_24, // @[:@131629.4]
  input  [63:0] io_ins_25, // @[:@131629.4]
  input  [63:0] io_ins_26, // @[:@131629.4]
  input  [63:0] io_ins_27, // @[:@131629.4]
  input  [63:0] io_ins_28, // @[:@131629.4]
  input  [63:0] io_ins_29, // @[:@131629.4]
  input  [63:0] io_ins_30, // @[:@131629.4]
  input  [63:0] io_ins_31, // @[:@131629.4]
  input  [63:0] io_ins_32, // @[:@131629.4]
  input  [63:0] io_ins_33, // @[:@131629.4]
  input  [63:0] io_ins_34, // @[:@131629.4]
  input  [63:0] io_ins_35, // @[:@131629.4]
  input  [63:0] io_ins_36, // @[:@131629.4]
  input  [63:0] io_ins_37, // @[:@131629.4]
  input  [63:0] io_ins_38, // @[:@131629.4]
  input  [63:0] io_ins_39, // @[:@131629.4]
  input  [63:0] io_ins_40, // @[:@131629.4]
  input  [63:0] io_ins_41, // @[:@131629.4]
  input  [63:0] io_ins_42, // @[:@131629.4]
  input  [63:0] io_ins_43, // @[:@131629.4]
  input  [63:0] io_ins_44, // @[:@131629.4]
  input  [63:0] io_ins_45, // @[:@131629.4]
  input  [63:0] io_ins_46, // @[:@131629.4]
  input  [63:0] io_ins_47, // @[:@131629.4]
  input  [63:0] io_ins_48, // @[:@131629.4]
  input  [63:0] io_ins_49, // @[:@131629.4]
  input  [63:0] io_ins_50, // @[:@131629.4]
  input  [63:0] io_ins_51, // @[:@131629.4]
  input  [63:0] io_ins_52, // @[:@131629.4]
  input  [63:0] io_ins_53, // @[:@131629.4]
  input  [63:0] io_ins_54, // @[:@131629.4]
  input  [63:0] io_ins_55, // @[:@131629.4]
  input  [63:0] io_ins_56, // @[:@131629.4]
  input  [63:0] io_ins_57, // @[:@131629.4]
  input  [63:0] io_ins_58, // @[:@131629.4]
  input  [63:0] io_ins_59, // @[:@131629.4]
  input  [63:0] io_ins_60, // @[:@131629.4]
  input  [63:0] io_ins_61, // @[:@131629.4]
  input  [63:0] io_ins_62, // @[:@131629.4]
  input  [63:0] io_ins_63, // @[:@131629.4]
  input  [63:0] io_ins_64, // @[:@131629.4]
  input  [63:0] io_ins_65, // @[:@131629.4]
  input  [63:0] io_ins_66, // @[:@131629.4]
  input  [63:0] io_ins_67, // @[:@131629.4]
  input  [63:0] io_ins_68, // @[:@131629.4]
  input  [63:0] io_ins_69, // @[:@131629.4]
  input  [63:0] io_ins_70, // @[:@131629.4]
  input  [63:0] io_ins_71, // @[:@131629.4]
  input  [63:0] io_ins_72, // @[:@131629.4]
  input  [63:0] io_ins_73, // @[:@131629.4]
  input  [63:0] io_ins_74, // @[:@131629.4]
  input  [63:0] io_ins_75, // @[:@131629.4]
  input  [63:0] io_ins_76, // @[:@131629.4]
  input  [63:0] io_ins_77, // @[:@131629.4]
  input  [63:0] io_ins_78, // @[:@131629.4]
  input  [63:0] io_ins_79, // @[:@131629.4]
  input  [63:0] io_ins_80, // @[:@131629.4]
  input  [63:0] io_ins_81, // @[:@131629.4]
  input  [63:0] io_ins_82, // @[:@131629.4]
  input  [63:0] io_ins_83, // @[:@131629.4]
  input  [63:0] io_ins_84, // @[:@131629.4]
  input  [63:0] io_ins_85, // @[:@131629.4]
  input  [63:0] io_ins_86, // @[:@131629.4]
  input  [63:0] io_ins_87, // @[:@131629.4]
  input  [63:0] io_ins_88, // @[:@131629.4]
  input  [63:0] io_ins_89, // @[:@131629.4]
  input  [63:0] io_ins_90, // @[:@131629.4]
  input  [63:0] io_ins_91, // @[:@131629.4]
  input  [63:0] io_ins_92, // @[:@131629.4]
  input  [63:0] io_ins_93, // @[:@131629.4]
  input  [63:0] io_ins_94, // @[:@131629.4]
  input  [63:0] io_ins_95, // @[:@131629.4]
  input  [63:0] io_ins_96, // @[:@131629.4]
  input  [63:0] io_ins_97, // @[:@131629.4]
  input  [63:0] io_ins_98, // @[:@131629.4]
  input  [63:0] io_ins_99, // @[:@131629.4]
  input  [63:0] io_ins_100, // @[:@131629.4]
  input  [63:0] io_ins_101, // @[:@131629.4]
  input  [63:0] io_ins_102, // @[:@131629.4]
  input  [63:0] io_ins_103, // @[:@131629.4]
  input  [63:0] io_ins_104, // @[:@131629.4]
  input  [63:0] io_ins_105, // @[:@131629.4]
  input  [63:0] io_ins_106, // @[:@131629.4]
  input  [63:0] io_ins_107, // @[:@131629.4]
  input  [63:0] io_ins_108, // @[:@131629.4]
  input  [63:0] io_ins_109, // @[:@131629.4]
  input  [63:0] io_ins_110, // @[:@131629.4]
  input  [63:0] io_ins_111, // @[:@131629.4]
  input  [63:0] io_ins_112, // @[:@131629.4]
  input  [63:0] io_ins_113, // @[:@131629.4]
  input  [63:0] io_ins_114, // @[:@131629.4]
  input  [63:0] io_ins_115, // @[:@131629.4]
  input  [63:0] io_ins_116, // @[:@131629.4]
  input  [63:0] io_ins_117, // @[:@131629.4]
  input  [63:0] io_ins_118, // @[:@131629.4]
  input  [63:0] io_ins_119, // @[:@131629.4]
  input  [63:0] io_ins_120, // @[:@131629.4]
  input  [63:0] io_ins_121, // @[:@131629.4]
  input  [63:0] io_ins_122, // @[:@131629.4]
  input  [63:0] io_ins_123, // @[:@131629.4]
  input  [63:0] io_ins_124, // @[:@131629.4]
  input  [63:0] io_ins_125, // @[:@131629.4]
  input  [63:0] io_ins_126, // @[:@131629.4]
  input  [63:0] io_ins_127, // @[:@131629.4]
  input  [63:0] io_ins_128, // @[:@131629.4]
  input  [63:0] io_ins_129, // @[:@131629.4]
  input  [63:0] io_ins_130, // @[:@131629.4]
  input  [63:0] io_ins_131, // @[:@131629.4]
  input  [63:0] io_ins_132, // @[:@131629.4]
  input  [63:0] io_ins_133, // @[:@131629.4]
  input  [63:0] io_ins_134, // @[:@131629.4]
  input  [63:0] io_ins_135, // @[:@131629.4]
  input  [63:0] io_ins_136, // @[:@131629.4]
  input  [63:0] io_ins_137, // @[:@131629.4]
  input  [63:0] io_ins_138, // @[:@131629.4]
  input  [63:0] io_ins_139, // @[:@131629.4]
  input  [63:0] io_ins_140, // @[:@131629.4]
  input  [63:0] io_ins_141, // @[:@131629.4]
  input  [63:0] io_ins_142, // @[:@131629.4]
  input  [63:0] io_ins_143, // @[:@131629.4]
  input  [63:0] io_ins_144, // @[:@131629.4]
  input  [63:0] io_ins_145, // @[:@131629.4]
  input  [63:0] io_ins_146, // @[:@131629.4]
  input  [63:0] io_ins_147, // @[:@131629.4]
  input  [63:0] io_ins_148, // @[:@131629.4]
  input  [63:0] io_ins_149, // @[:@131629.4]
  input  [63:0] io_ins_150, // @[:@131629.4]
  input  [63:0] io_ins_151, // @[:@131629.4]
  input  [63:0] io_ins_152, // @[:@131629.4]
  input  [63:0] io_ins_153, // @[:@131629.4]
  input  [63:0] io_ins_154, // @[:@131629.4]
  input  [63:0] io_ins_155, // @[:@131629.4]
  input  [63:0] io_ins_156, // @[:@131629.4]
  input  [63:0] io_ins_157, // @[:@131629.4]
  input  [63:0] io_ins_158, // @[:@131629.4]
  input  [63:0] io_ins_159, // @[:@131629.4]
  input  [63:0] io_ins_160, // @[:@131629.4]
  input  [63:0] io_ins_161, // @[:@131629.4]
  input  [63:0] io_ins_162, // @[:@131629.4]
  input  [63:0] io_ins_163, // @[:@131629.4]
  input  [63:0] io_ins_164, // @[:@131629.4]
  input  [63:0] io_ins_165, // @[:@131629.4]
  input  [63:0] io_ins_166, // @[:@131629.4]
  input  [63:0] io_ins_167, // @[:@131629.4]
  input  [63:0] io_ins_168, // @[:@131629.4]
  input  [63:0] io_ins_169, // @[:@131629.4]
  input  [63:0] io_ins_170, // @[:@131629.4]
  input  [63:0] io_ins_171, // @[:@131629.4]
  input  [63:0] io_ins_172, // @[:@131629.4]
  input  [63:0] io_ins_173, // @[:@131629.4]
  input  [63:0] io_ins_174, // @[:@131629.4]
  input  [63:0] io_ins_175, // @[:@131629.4]
  input  [63:0] io_ins_176, // @[:@131629.4]
  input  [63:0] io_ins_177, // @[:@131629.4]
  input  [63:0] io_ins_178, // @[:@131629.4]
  input  [63:0] io_ins_179, // @[:@131629.4]
  input  [63:0] io_ins_180, // @[:@131629.4]
  input  [63:0] io_ins_181, // @[:@131629.4]
  input  [63:0] io_ins_182, // @[:@131629.4]
  input  [63:0] io_ins_183, // @[:@131629.4]
  input  [63:0] io_ins_184, // @[:@131629.4]
  input  [63:0] io_ins_185, // @[:@131629.4]
  input  [63:0] io_ins_186, // @[:@131629.4]
  input  [63:0] io_ins_187, // @[:@131629.4]
  input  [63:0] io_ins_188, // @[:@131629.4]
  input  [63:0] io_ins_189, // @[:@131629.4]
  input  [63:0] io_ins_190, // @[:@131629.4]
  input  [63:0] io_ins_191, // @[:@131629.4]
  input  [63:0] io_ins_192, // @[:@131629.4]
  input  [63:0] io_ins_193, // @[:@131629.4]
  input  [63:0] io_ins_194, // @[:@131629.4]
  input  [63:0] io_ins_195, // @[:@131629.4]
  input  [63:0] io_ins_196, // @[:@131629.4]
  input  [63:0] io_ins_197, // @[:@131629.4]
  input  [63:0] io_ins_198, // @[:@131629.4]
  input  [63:0] io_ins_199, // @[:@131629.4]
  input  [63:0] io_ins_200, // @[:@131629.4]
  input  [63:0] io_ins_201, // @[:@131629.4]
  input  [63:0] io_ins_202, // @[:@131629.4]
  input  [63:0] io_ins_203, // @[:@131629.4]
  input  [63:0] io_ins_204, // @[:@131629.4]
  input  [63:0] io_ins_205, // @[:@131629.4]
  input  [63:0] io_ins_206, // @[:@131629.4]
  input  [63:0] io_ins_207, // @[:@131629.4]
  input  [63:0] io_ins_208, // @[:@131629.4]
  input  [63:0] io_ins_209, // @[:@131629.4]
  input  [63:0] io_ins_210, // @[:@131629.4]
  input  [63:0] io_ins_211, // @[:@131629.4]
  input  [63:0] io_ins_212, // @[:@131629.4]
  input  [63:0] io_ins_213, // @[:@131629.4]
  input  [63:0] io_ins_214, // @[:@131629.4]
  input  [63:0] io_ins_215, // @[:@131629.4]
  input  [63:0] io_ins_216, // @[:@131629.4]
  input  [63:0] io_ins_217, // @[:@131629.4]
  input  [63:0] io_ins_218, // @[:@131629.4]
  input  [63:0] io_ins_219, // @[:@131629.4]
  input  [63:0] io_ins_220, // @[:@131629.4]
  input  [63:0] io_ins_221, // @[:@131629.4]
  input  [63:0] io_ins_222, // @[:@131629.4]
  input  [63:0] io_ins_223, // @[:@131629.4]
  input  [63:0] io_ins_224, // @[:@131629.4]
  input  [63:0] io_ins_225, // @[:@131629.4]
  input  [63:0] io_ins_226, // @[:@131629.4]
  input  [63:0] io_ins_227, // @[:@131629.4]
  input  [63:0] io_ins_228, // @[:@131629.4]
  input  [63:0] io_ins_229, // @[:@131629.4]
  input  [63:0] io_ins_230, // @[:@131629.4]
  input  [63:0] io_ins_231, // @[:@131629.4]
  input  [63:0] io_ins_232, // @[:@131629.4]
  input  [63:0] io_ins_233, // @[:@131629.4]
  input  [63:0] io_ins_234, // @[:@131629.4]
  input  [63:0] io_ins_235, // @[:@131629.4]
  input  [63:0] io_ins_236, // @[:@131629.4]
  input  [63:0] io_ins_237, // @[:@131629.4]
  input  [63:0] io_ins_238, // @[:@131629.4]
  input  [63:0] io_ins_239, // @[:@131629.4]
  input  [63:0] io_ins_240, // @[:@131629.4]
  input  [63:0] io_ins_241, // @[:@131629.4]
  input  [63:0] io_ins_242, // @[:@131629.4]
  input  [63:0] io_ins_243, // @[:@131629.4]
  input  [63:0] io_ins_244, // @[:@131629.4]
  input  [63:0] io_ins_245, // @[:@131629.4]
  input  [63:0] io_ins_246, // @[:@131629.4]
  input  [63:0] io_ins_247, // @[:@131629.4]
  input  [63:0] io_ins_248, // @[:@131629.4]
  input  [63:0] io_ins_249, // @[:@131629.4]
  input  [63:0] io_ins_250, // @[:@131629.4]
  input  [63:0] io_ins_251, // @[:@131629.4]
  input  [63:0] io_ins_252, // @[:@131629.4]
  input  [63:0] io_ins_253, // @[:@131629.4]
  input  [63:0] io_ins_254, // @[:@131629.4]
  input  [63:0] io_ins_255, // @[:@131629.4]
  input  [63:0] io_ins_256, // @[:@131629.4]
  input  [63:0] io_ins_257, // @[:@131629.4]
  input  [63:0] io_ins_258, // @[:@131629.4]
  input  [63:0] io_ins_259, // @[:@131629.4]
  input  [63:0] io_ins_260, // @[:@131629.4]
  input  [63:0] io_ins_261, // @[:@131629.4]
  input  [63:0] io_ins_262, // @[:@131629.4]
  input  [63:0] io_ins_263, // @[:@131629.4]
  input  [63:0] io_ins_264, // @[:@131629.4]
  input  [63:0] io_ins_265, // @[:@131629.4]
  input  [63:0] io_ins_266, // @[:@131629.4]
  input  [63:0] io_ins_267, // @[:@131629.4]
  input  [63:0] io_ins_268, // @[:@131629.4]
  input  [63:0] io_ins_269, // @[:@131629.4]
  input  [63:0] io_ins_270, // @[:@131629.4]
  input  [63:0] io_ins_271, // @[:@131629.4]
  input  [63:0] io_ins_272, // @[:@131629.4]
  input  [63:0] io_ins_273, // @[:@131629.4]
  input  [63:0] io_ins_274, // @[:@131629.4]
  input  [63:0] io_ins_275, // @[:@131629.4]
  input  [63:0] io_ins_276, // @[:@131629.4]
  input  [63:0] io_ins_277, // @[:@131629.4]
  input  [63:0] io_ins_278, // @[:@131629.4]
  input  [63:0] io_ins_279, // @[:@131629.4]
  input  [63:0] io_ins_280, // @[:@131629.4]
  input  [63:0] io_ins_281, // @[:@131629.4]
  input  [63:0] io_ins_282, // @[:@131629.4]
  input  [63:0] io_ins_283, // @[:@131629.4]
  input  [63:0] io_ins_284, // @[:@131629.4]
  input  [63:0] io_ins_285, // @[:@131629.4]
  input  [63:0] io_ins_286, // @[:@131629.4]
  input  [63:0] io_ins_287, // @[:@131629.4]
  input  [63:0] io_ins_288, // @[:@131629.4]
  input  [63:0] io_ins_289, // @[:@131629.4]
  input  [63:0] io_ins_290, // @[:@131629.4]
  input  [63:0] io_ins_291, // @[:@131629.4]
  input  [63:0] io_ins_292, // @[:@131629.4]
  input  [63:0] io_ins_293, // @[:@131629.4]
  input  [63:0] io_ins_294, // @[:@131629.4]
  input  [63:0] io_ins_295, // @[:@131629.4]
  input  [63:0] io_ins_296, // @[:@131629.4]
  input  [63:0] io_ins_297, // @[:@131629.4]
  input  [63:0] io_ins_298, // @[:@131629.4]
  input  [63:0] io_ins_299, // @[:@131629.4]
  input  [63:0] io_ins_300, // @[:@131629.4]
  input  [63:0] io_ins_301, // @[:@131629.4]
  input  [63:0] io_ins_302, // @[:@131629.4]
  input  [63:0] io_ins_303, // @[:@131629.4]
  input  [63:0] io_ins_304, // @[:@131629.4]
  input  [63:0] io_ins_305, // @[:@131629.4]
  input  [63:0] io_ins_306, // @[:@131629.4]
  input  [63:0] io_ins_307, // @[:@131629.4]
  input  [63:0] io_ins_308, // @[:@131629.4]
  input  [63:0] io_ins_309, // @[:@131629.4]
  input  [63:0] io_ins_310, // @[:@131629.4]
  input  [63:0] io_ins_311, // @[:@131629.4]
  input  [63:0] io_ins_312, // @[:@131629.4]
  input  [63:0] io_ins_313, // @[:@131629.4]
  input  [63:0] io_ins_314, // @[:@131629.4]
  input  [63:0] io_ins_315, // @[:@131629.4]
  input  [63:0] io_ins_316, // @[:@131629.4]
  input  [63:0] io_ins_317, // @[:@131629.4]
  input  [63:0] io_ins_318, // @[:@131629.4]
  input  [63:0] io_ins_319, // @[:@131629.4]
  input  [63:0] io_ins_320, // @[:@131629.4]
  input  [63:0] io_ins_321, // @[:@131629.4]
  input  [63:0] io_ins_322, // @[:@131629.4]
  input  [63:0] io_ins_323, // @[:@131629.4]
  input  [63:0] io_ins_324, // @[:@131629.4]
  input  [63:0] io_ins_325, // @[:@131629.4]
  input  [63:0] io_ins_326, // @[:@131629.4]
  input  [63:0] io_ins_327, // @[:@131629.4]
  input  [63:0] io_ins_328, // @[:@131629.4]
  input  [63:0] io_ins_329, // @[:@131629.4]
  input  [63:0] io_ins_330, // @[:@131629.4]
  input  [63:0] io_ins_331, // @[:@131629.4]
  input  [63:0] io_ins_332, // @[:@131629.4]
  input  [63:0] io_ins_333, // @[:@131629.4]
  input  [63:0] io_ins_334, // @[:@131629.4]
  input  [63:0] io_ins_335, // @[:@131629.4]
  input  [63:0] io_ins_336, // @[:@131629.4]
  input  [63:0] io_ins_337, // @[:@131629.4]
  input  [63:0] io_ins_338, // @[:@131629.4]
  input  [63:0] io_ins_339, // @[:@131629.4]
  input  [63:0] io_ins_340, // @[:@131629.4]
  input  [63:0] io_ins_341, // @[:@131629.4]
  input  [63:0] io_ins_342, // @[:@131629.4]
  input  [63:0] io_ins_343, // @[:@131629.4]
  input  [63:0] io_ins_344, // @[:@131629.4]
  input  [63:0] io_ins_345, // @[:@131629.4]
  input  [63:0] io_ins_346, // @[:@131629.4]
  input  [63:0] io_ins_347, // @[:@131629.4]
  input  [63:0] io_ins_348, // @[:@131629.4]
  input  [63:0] io_ins_349, // @[:@131629.4]
  input  [63:0] io_ins_350, // @[:@131629.4]
  input  [63:0] io_ins_351, // @[:@131629.4]
  input  [63:0] io_ins_352, // @[:@131629.4]
  input  [63:0] io_ins_353, // @[:@131629.4]
  input  [63:0] io_ins_354, // @[:@131629.4]
  input  [63:0] io_ins_355, // @[:@131629.4]
  input  [63:0] io_ins_356, // @[:@131629.4]
  input  [63:0] io_ins_357, // @[:@131629.4]
  input  [63:0] io_ins_358, // @[:@131629.4]
  input  [63:0] io_ins_359, // @[:@131629.4]
  input  [63:0] io_ins_360, // @[:@131629.4]
  input  [63:0] io_ins_361, // @[:@131629.4]
  input  [63:0] io_ins_362, // @[:@131629.4]
  input  [63:0] io_ins_363, // @[:@131629.4]
  input  [63:0] io_ins_364, // @[:@131629.4]
  input  [63:0] io_ins_365, // @[:@131629.4]
  input  [63:0] io_ins_366, // @[:@131629.4]
  input  [63:0] io_ins_367, // @[:@131629.4]
  input  [63:0] io_ins_368, // @[:@131629.4]
  input  [63:0] io_ins_369, // @[:@131629.4]
  input  [63:0] io_ins_370, // @[:@131629.4]
  input  [63:0] io_ins_371, // @[:@131629.4]
  input  [63:0] io_ins_372, // @[:@131629.4]
  input  [63:0] io_ins_373, // @[:@131629.4]
  input  [63:0] io_ins_374, // @[:@131629.4]
  input  [63:0] io_ins_375, // @[:@131629.4]
  input  [63:0] io_ins_376, // @[:@131629.4]
  input  [63:0] io_ins_377, // @[:@131629.4]
  input  [63:0] io_ins_378, // @[:@131629.4]
  input  [63:0] io_ins_379, // @[:@131629.4]
  input  [63:0] io_ins_380, // @[:@131629.4]
  input  [63:0] io_ins_381, // @[:@131629.4]
  input  [63:0] io_ins_382, // @[:@131629.4]
  input  [63:0] io_ins_383, // @[:@131629.4]
  input  [63:0] io_ins_384, // @[:@131629.4]
  input  [63:0] io_ins_385, // @[:@131629.4]
  input  [63:0] io_ins_386, // @[:@131629.4]
  input  [63:0] io_ins_387, // @[:@131629.4]
  input  [63:0] io_ins_388, // @[:@131629.4]
  input  [63:0] io_ins_389, // @[:@131629.4]
  input  [63:0] io_ins_390, // @[:@131629.4]
  input  [63:0] io_ins_391, // @[:@131629.4]
  input  [63:0] io_ins_392, // @[:@131629.4]
  input  [63:0] io_ins_393, // @[:@131629.4]
  input  [63:0] io_ins_394, // @[:@131629.4]
  input  [63:0] io_ins_395, // @[:@131629.4]
  input  [63:0] io_ins_396, // @[:@131629.4]
  input  [63:0] io_ins_397, // @[:@131629.4]
  input  [63:0] io_ins_398, // @[:@131629.4]
  input  [63:0] io_ins_399, // @[:@131629.4]
  input  [63:0] io_ins_400, // @[:@131629.4]
  input  [63:0] io_ins_401, // @[:@131629.4]
  input  [63:0] io_ins_402, // @[:@131629.4]
  input  [63:0] io_ins_403, // @[:@131629.4]
  input  [63:0] io_ins_404, // @[:@131629.4]
  input  [63:0] io_ins_405, // @[:@131629.4]
  input  [63:0] io_ins_406, // @[:@131629.4]
  input  [63:0] io_ins_407, // @[:@131629.4]
  input  [63:0] io_ins_408, // @[:@131629.4]
  input  [63:0] io_ins_409, // @[:@131629.4]
  input  [63:0] io_ins_410, // @[:@131629.4]
  input  [63:0] io_ins_411, // @[:@131629.4]
  input  [63:0] io_ins_412, // @[:@131629.4]
  input  [63:0] io_ins_413, // @[:@131629.4]
  input  [63:0] io_ins_414, // @[:@131629.4]
  input  [63:0] io_ins_415, // @[:@131629.4]
  input  [63:0] io_ins_416, // @[:@131629.4]
  input  [63:0] io_ins_417, // @[:@131629.4]
  input  [63:0] io_ins_418, // @[:@131629.4]
  input  [63:0] io_ins_419, // @[:@131629.4]
  input  [63:0] io_ins_420, // @[:@131629.4]
  input  [63:0] io_ins_421, // @[:@131629.4]
  input  [63:0] io_ins_422, // @[:@131629.4]
  input  [63:0] io_ins_423, // @[:@131629.4]
  input  [63:0] io_ins_424, // @[:@131629.4]
  input  [63:0] io_ins_425, // @[:@131629.4]
  input  [63:0] io_ins_426, // @[:@131629.4]
  input  [63:0] io_ins_427, // @[:@131629.4]
  input  [63:0] io_ins_428, // @[:@131629.4]
  input  [63:0] io_ins_429, // @[:@131629.4]
  input  [63:0] io_ins_430, // @[:@131629.4]
  input  [63:0] io_ins_431, // @[:@131629.4]
  input  [63:0] io_ins_432, // @[:@131629.4]
  input  [63:0] io_ins_433, // @[:@131629.4]
  input  [63:0] io_ins_434, // @[:@131629.4]
  input  [63:0] io_ins_435, // @[:@131629.4]
  input  [63:0] io_ins_436, // @[:@131629.4]
  input  [63:0] io_ins_437, // @[:@131629.4]
  input  [63:0] io_ins_438, // @[:@131629.4]
  input  [63:0] io_ins_439, // @[:@131629.4]
  input  [63:0] io_ins_440, // @[:@131629.4]
  input  [63:0] io_ins_441, // @[:@131629.4]
  input  [63:0] io_ins_442, // @[:@131629.4]
  input  [63:0] io_ins_443, // @[:@131629.4]
  input  [63:0] io_ins_444, // @[:@131629.4]
  input  [63:0] io_ins_445, // @[:@131629.4]
  input  [63:0] io_ins_446, // @[:@131629.4]
  input  [63:0] io_ins_447, // @[:@131629.4]
  input  [63:0] io_ins_448, // @[:@131629.4]
  input  [63:0] io_ins_449, // @[:@131629.4]
  input  [63:0] io_ins_450, // @[:@131629.4]
  input  [63:0] io_ins_451, // @[:@131629.4]
  input  [63:0] io_ins_452, // @[:@131629.4]
  input  [63:0] io_ins_453, // @[:@131629.4]
  input  [63:0] io_ins_454, // @[:@131629.4]
  input  [63:0] io_ins_455, // @[:@131629.4]
  input  [63:0] io_ins_456, // @[:@131629.4]
  input  [63:0] io_ins_457, // @[:@131629.4]
  input  [63:0] io_ins_458, // @[:@131629.4]
  input  [63:0] io_ins_459, // @[:@131629.4]
  input  [63:0] io_ins_460, // @[:@131629.4]
  input  [63:0] io_ins_461, // @[:@131629.4]
  input  [63:0] io_ins_462, // @[:@131629.4]
  input  [63:0] io_ins_463, // @[:@131629.4]
  input  [63:0] io_ins_464, // @[:@131629.4]
  input  [63:0] io_ins_465, // @[:@131629.4]
  input  [63:0] io_ins_466, // @[:@131629.4]
  input  [63:0] io_ins_467, // @[:@131629.4]
  input  [63:0] io_ins_468, // @[:@131629.4]
  input  [63:0] io_ins_469, // @[:@131629.4]
  input  [63:0] io_ins_470, // @[:@131629.4]
  input  [63:0] io_ins_471, // @[:@131629.4]
  input  [63:0] io_ins_472, // @[:@131629.4]
  input  [63:0] io_ins_473, // @[:@131629.4]
  input  [63:0] io_ins_474, // @[:@131629.4]
  input  [63:0] io_ins_475, // @[:@131629.4]
  input  [63:0] io_ins_476, // @[:@131629.4]
  input  [63:0] io_ins_477, // @[:@131629.4]
  input  [63:0] io_ins_478, // @[:@131629.4]
  input  [63:0] io_ins_479, // @[:@131629.4]
  input  [63:0] io_ins_480, // @[:@131629.4]
  input  [63:0] io_ins_481, // @[:@131629.4]
  input  [63:0] io_ins_482, // @[:@131629.4]
  input  [63:0] io_ins_483, // @[:@131629.4]
  input  [63:0] io_ins_484, // @[:@131629.4]
  input  [63:0] io_ins_485, // @[:@131629.4]
  input  [63:0] io_ins_486, // @[:@131629.4]
  input  [63:0] io_ins_487, // @[:@131629.4]
  input  [63:0] io_ins_488, // @[:@131629.4]
  input  [63:0] io_ins_489, // @[:@131629.4]
  input  [63:0] io_ins_490, // @[:@131629.4]
  input  [63:0] io_ins_491, // @[:@131629.4]
  input  [63:0] io_ins_492, // @[:@131629.4]
  input  [63:0] io_ins_493, // @[:@131629.4]
  input  [63:0] io_ins_494, // @[:@131629.4]
  input  [63:0] io_ins_495, // @[:@131629.4]
  input  [63:0] io_ins_496, // @[:@131629.4]
  input  [63:0] io_ins_497, // @[:@131629.4]
  input  [63:0] io_ins_498, // @[:@131629.4]
  input  [63:0] io_ins_499, // @[:@131629.4]
  input  [63:0] io_ins_500, // @[:@131629.4]
  input  [63:0] io_ins_501, // @[:@131629.4]
  input  [63:0] io_ins_502, // @[:@131629.4]
  input  [8:0]  io_sel, // @[:@131629.4]
  output [63:0] io_out // @[:@131629.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@131631.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@131631.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@131631.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@131631.4]
endmodule
module RegFile( // @[:@131633.2]
  input         clock, // @[:@131634.4]
  input         reset, // @[:@131635.4]
  input  [31:0] io_raddr, // @[:@131636.4]
  input         io_wen, // @[:@131636.4]
  input  [31:0] io_waddr, // @[:@131636.4]
  input  [63:0] io_wdata, // @[:@131636.4]
  output [63:0] io_rdata, // @[:@131636.4]
  input         io_reset, // @[:@131636.4]
  output [63:0] io_argIns_0, // @[:@131636.4]
  output [63:0] io_argIns_1, // @[:@131636.4]
  output [63:0] io_argIns_2, // @[:@131636.4]
  output [63:0] io_argIns_3, // @[:@131636.4]
  input         io_argOuts_0_valid, // @[:@131636.4]
  input  [63:0] io_argOuts_0_bits, // @[:@131636.4]
  input         io_argOuts_1_valid, // @[:@131636.4]
  input  [63:0] io_argOuts_1_bits // @[:@131636.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@133646.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@133646.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@133646.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@133658.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@133658.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@133658.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@133658.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@133658.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@133658.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@133677.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@133677.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@133677.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@133677.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@133677.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@133677.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@133689.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@133689.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@133701.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@133701.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@133701.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@133701.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@133701.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@133701.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@133715.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@133715.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@133715.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@133715.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@133715.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@133715.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@133729.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@133729.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@133729.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@133729.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@133729.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@133729.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@133743.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@133743.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@133743.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@133743.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@133743.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@133743.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@133757.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@133757.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@133757.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@133757.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@133757.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@133757.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@133771.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@133771.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@133771.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@133771.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@133771.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@133771.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@133785.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@133785.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@133785.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@133785.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@133785.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@133785.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@133799.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@133799.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@133799.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@133799.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@133799.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@133799.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@133813.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@133813.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@133813.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@133813.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@133813.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@133813.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@133827.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@133827.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@133827.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@133827.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@133827.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@133827.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@133841.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@133841.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@133841.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@133841.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@133841.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@133841.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@133855.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@133855.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@133855.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@133855.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@133855.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@133855.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@133869.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@133869.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@133869.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@133869.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@133869.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@133869.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@133883.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@133883.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@133883.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@133883.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@133883.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@133883.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@133897.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@133897.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@133897.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@133897.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@133897.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@133897.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@133911.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@133911.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@133911.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@133911.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@133911.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@133911.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@133925.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@133925.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@133925.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@133925.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@133925.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@133925.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@133939.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@133939.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@133939.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@133939.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@133939.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@133939.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@133953.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@133953.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@133953.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@133953.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@133953.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@133953.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@133967.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@133967.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@133967.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@133967.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@133967.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@133967.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@133981.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@133981.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@133981.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@133981.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@133981.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@133981.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@133995.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@133995.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@133995.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@133995.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@133995.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@133995.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@134009.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@134009.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@134009.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@134009.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@134009.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@134009.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@134023.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@134023.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@134023.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@134023.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@134023.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@134023.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@134037.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@134037.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@134037.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@134037.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@134037.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@134037.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@134051.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@134051.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@134051.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@134051.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@134051.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@134051.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@134065.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@134065.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@134065.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@134065.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@134065.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@134065.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@134079.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@134079.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@134079.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@134079.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@134079.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@134079.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@134093.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@134093.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@134093.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@134093.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@134093.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@134093.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@134107.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@134107.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@134107.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@134107.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@134107.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@134107.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@134121.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@134121.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@134121.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@134121.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@134121.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@134121.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@134135.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@134135.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@134135.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@134135.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@134135.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@134135.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@134149.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@134149.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@134149.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@134149.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@134149.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@134149.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@134163.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@134163.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@134163.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@134163.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@134163.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@134163.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@134177.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@134177.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@134177.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@134177.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@134177.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@134177.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@134191.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@134191.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@134191.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@134191.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@134191.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@134191.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@134205.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@134205.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@134205.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@134205.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@134205.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@134205.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@134219.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@134219.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@134219.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@134219.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@134219.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@134219.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@134233.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@134233.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@134233.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@134233.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@134233.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@134233.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@134247.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@134247.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@134247.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@134247.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@134247.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@134247.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@134261.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@134261.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@134261.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@134261.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@134261.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@134261.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@134275.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@134275.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@134275.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@134275.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@134275.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@134275.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@134289.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@134289.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@134289.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@134289.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@134289.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@134289.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@134303.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@134303.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@134303.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@134303.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@134303.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@134303.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@134317.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@134317.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@134317.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@134317.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@134317.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@134317.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@134331.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@134331.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@134331.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@134331.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@134331.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@134331.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@134345.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@134345.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@134345.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@134345.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@134345.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@134345.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@134359.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@134359.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@134359.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@134359.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@134359.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@134359.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@134373.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@134373.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@134373.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@134373.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@134373.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@134373.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@134387.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@134387.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@134387.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@134387.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@134387.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@134387.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@134401.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@134401.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@134401.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@134401.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@134401.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@134401.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@134415.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@134415.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@134415.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@134415.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@134415.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@134415.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@134429.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@134429.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@134429.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@134429.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@134429.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@134429.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@134443.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@134443.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@134443.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@134443.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@134443.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@134443.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@134457.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@134457.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@134457.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@134457.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@134457.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@134457.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@134471.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@134471.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@134471.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@134471.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@134471.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@134471.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@134485.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@134485.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@134485.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@134485.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@134485.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@134485.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@134499.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@134499.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@134499.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@134499.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@134499.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@134499.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@134513.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@134513.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@134513.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@134513.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@134513.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@134513.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@134527.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@134527.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@134527.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@134527.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@134527.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@134527.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@134541.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@134541.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@134541.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@134541.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@134541.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@134541.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@134555.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@134555.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@134555.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@134555.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@134555.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@134555.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@134569.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@134569.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@134569.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@134569.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@134569.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@134569.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@134583.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@134583.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@134583.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@134583.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@134583.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@134583.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@134597.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@134597.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@134597.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@134597.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@134597.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@134597.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@134611.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@134611.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@134611.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@134611.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@134611.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@134611.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@134625.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@134625.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@134625.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@134625.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@134625.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@134625.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@134639.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@134639.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@134639.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@134639.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@134639.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@134639.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@134653.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@134653.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@134653.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@134653.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@134653.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@134653.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@134667.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@134667.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@134667.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@134667.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@134667.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@134667.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@134681.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@134681.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@134681.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@134681.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@134681.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@134681.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@134695.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@134695.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@134695.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@134695.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@134695.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@134695.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@134709.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@134709.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@134709.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@134709.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@134709.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@134709.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@134723.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@134723.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@134723.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@134723.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@134723.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@134723.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@134737.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@134737.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@134737.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@134737.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@134737.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@134737.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@134751.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@134751.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@134751.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@134751.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@134751.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@134751.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@134765.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@134765.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@134765.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@134765.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@134765.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@134765.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@134779.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@134779.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@134779.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@134779.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@134779.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@134779.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@134793.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@134793.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@134793.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@134793.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@134793.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@134793.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@134807.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@134807.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@134807.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@134807.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@134807.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@134807.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@134821.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@134821.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@134821.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@134821.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@134821.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@134821.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@134835.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@134835.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@134835.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@134835.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@134835.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@134835.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@134849.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@134849.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@134849.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@134849.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@134849.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@134849.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@134863.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@134863.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@134863.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@134863.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@134863.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@134863.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@134877.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@134877.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@134877.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@134877.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@134877.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@134877.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@134891.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@134891.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@134891.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@134891.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@134891.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@134891.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@134905.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@134905.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@134905.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@134905.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@134905.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@134905.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@134919.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@134919.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@134919.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@134919.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@134919.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@134919.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@134933.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@134933.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@134933.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@134933.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@134933.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@134933.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@134947.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@134947.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@134947.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@134947.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@134947.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@134947.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@134961.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@134961.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@134961.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@134961.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@134961.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@134961.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@134975.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@134975.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@134975.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@134975.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@134975.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@134975.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@134989.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@134989.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@134989.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@134989.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@134989.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@134989.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@135003.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@135003.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@135003.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@135003.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@135003.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@135003.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@135017.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@135017.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@135017.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@135017.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@135017.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@135017.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@135031.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@135031.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@135031.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@135031.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@135031.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@135031.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@135045.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@135045.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@135045.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@135045.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@135045.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@135045.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@135059.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@135059.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@135059.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@135059.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@135059.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@135059.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@135073.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@135073.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@135073.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@135073.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@135073.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@135073.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@135087.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@135087.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@135087.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@135087.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@135087.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@135087.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@135101.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@135101.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@135101.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@135101.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@135101.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@135101.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@135115.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@135115.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@135115.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@135115.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@135115.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@135115.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@135129.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@135129.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@135129.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@135129.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@135129.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@135129.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@135143.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@135143.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@135143.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@135143.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@135143.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@135143.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@135157.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@135157.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@135157.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@135157.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@135157.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@135157.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@135171.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@135171.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@135171.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@135171.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@135171.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@135171.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@135185.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@135185.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@135185.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@135185.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@135185.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@135185.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@135199.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@135199.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@135199.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@135199.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@135199.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@135199.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@135213.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@135213.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@135213.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@135213.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@135213.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@135213.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@135227.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@135227.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@135227.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@135227.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@135227.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@135227.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@135241.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@135241.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@135241.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@135241.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@135241.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@135241.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@135255.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@135255.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@135255.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@135255.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@135255.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@135255.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@135269.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@135269.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@135269.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@135269.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@135269.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@135269.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@135283.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@135283.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@135283.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@135283.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@135283.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@135283.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@135297.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@135297.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@135297.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@135297.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@135297.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@135297.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@135311.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@135311.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@135311.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@135311.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@135311.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@135311.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@135325.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@135325.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@135325.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@135325.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@135325.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@135325.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@135339.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@135339.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@135339.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@135339.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@135339.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@135339.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@135353.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@135353.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@135353.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@135353.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@135353.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@135353.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@135367.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@135367.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@135367.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@135367.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@135367.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@135367.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@135381.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@135381.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@135381.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@135381.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@135381.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@135381.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@135395.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@135395.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@135395.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@135395.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@135395.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@135395.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@135409.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@135409.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@135409.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@135409.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@135409.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@135409.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@135423.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@135423.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@135423.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@135423.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@135423.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@135423.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@135437.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@135437.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@135437.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@135437.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@135437.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@135437.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@135451.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@135451.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@135451.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@135451.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@135451.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@135451.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@135465.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@135465.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@135465.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@135465.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@135465.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@135465.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@135479.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@135479.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@135479.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@135479.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@135479.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@135479.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@135493.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@135493.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@135493.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@135493.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@135493.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@135493.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@135507.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@135507.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@135507.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@135507.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@135507.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@135507.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@135521.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@135521.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@135521.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@135521.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@135521.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@135521.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@135535.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@135535.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@135535.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@135535.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@135535.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@135535.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@135549.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@135549.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@135549.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@135549.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@135549.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@135549.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@135563.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@135563.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@135563.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@135563.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@135563.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@135563.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@135577.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@135577.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@135577.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@135577.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@135577.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@135577.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@135591.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@135591.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@135591.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@135591.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@135591.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@135591.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@135605.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@135605.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@135605.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@135605.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@135605.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@135605.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@135619.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@135619.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@135619.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@135619.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@135619.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@135619.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@135633.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@135633.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@135633.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@135633.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@135633.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@135633.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@135647.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@135647.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@135647.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@135647.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@135647.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@135647.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@135661.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@135661.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@135661.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@135661.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@135661.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@135661.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@135675.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@135675.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@135675.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@135675.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@135675.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@135675.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@135689.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@135689.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@135689.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@135689.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@135689.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@135689.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@135703.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@135703.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@135703.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@135703.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@135703.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@135703.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@135717.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@135717.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@135717.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@135717.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@135717.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@135717.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@135731.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@135731.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@135731.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@135731.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@135731.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@135731.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@135745.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@135745.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@135745.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@135745.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@135745.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@135745.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@135759.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@135759.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@135759.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@135759.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@135759.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@135759.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@135773.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@135773.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@135773.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@135773.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@135773.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@135773.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@135787.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@135787.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@135787.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@135787.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@135787.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@135787.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@135801.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@135801.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@135801.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@135801.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@135801.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@135801.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@135815.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@135815.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@135815.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@135815.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@135815.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@135815.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@135829.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@135829.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@135829.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@135829.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@135829.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@135829.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@135843.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@135843.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@135843.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@135843.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@135843.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@135843.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@135857.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@135857.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@135857.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@135857.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@135857.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@135857.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@135871.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@135871.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@135871.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@135871.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@135871.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@135871.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@135885.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@135885.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@135885.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@135885.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@135885.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@135885.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@135899.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@135899.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@135899.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@135899.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@135899.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@135899.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@135913.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@135913.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@135913.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@135913.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@135913.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@135913.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@135927.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@135927.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@135927.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@135927.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@135927.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@135927.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@135941.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@135941.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@135941.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@135941.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@135941.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@135941.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@135955.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@135955.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@135955.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@135955.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@135955.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@135955.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@135969.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@135969.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@135969.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@135969.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@135969.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@135969.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@135983.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@135983.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@135983.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@135983.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@135983.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@135983.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@135997.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@135997.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@135997.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@135997.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@135997.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@135997.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@136011.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@136011.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@136011.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@136011.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@136011.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@136011.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@136025.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@136025.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@136025.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@136025.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@136025.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@136025.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@136039.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@136039.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@136039.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@136039.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@136039.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@136039.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@136053.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@136053.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@136053.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@136053.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@136053.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@136053.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@136067.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@136067.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@136067.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@136067.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@136067.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@136067.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@136081.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@136081.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@136081.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@136081.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@136081.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@136081.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@136095.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@136095.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@136095.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@136095.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@136095.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@136095.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@136109.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@136109.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@136109.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@136109.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@136109.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@136109.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@136123.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@136123.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@136123.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@136123.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@136123.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@136123.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@136137.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@136137.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@136137.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@136137.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@136137.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@136137.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@136151.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@136151.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@136151.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@136151.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@136151.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@136151.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@136165.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@136165.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@136165.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@136165.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@136165.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@136165.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@136179.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@136179.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@136179.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@136179.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@136179.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@136179.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@136193.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@136193.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@136193.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@136193.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@136193.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@136193.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@136207.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@136207.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@136207.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@136207.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@136207.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@136207.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@136221.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@136221.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@136221.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@136221.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@136221.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@136221.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@136235.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@136235.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@136235.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@136235.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@136235.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@136235.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@136249.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@136249.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@136249.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@136249.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@136249.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@136249.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@136263.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@136263.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@136263.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@136263.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@136263.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@136263.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@136277.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@136277.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@136277.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@136277.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@136277.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@136277.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@136291.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@136291.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@136291.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@136291.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@136291.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@136291.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@136305.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@136305.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@136305.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@136305.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@136305.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@136305.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@136319.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@136319.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@136319.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@136319.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@136319.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@136319.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@136333.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@136333.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@136333.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@136333.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@136333.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@136333.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@136347.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@136347.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@136347.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@136347.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@136347.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@136347.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@136361.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@136361.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@136361.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@136361.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@136361.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@136361.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@136375.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@136375.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@136375.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@136375.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@136375.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@136375.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@136389.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@136389.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@136389.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@136389.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@136389.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@136389.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@136403.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@136403.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@136403.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@136403.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@136403.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@136403.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@136417.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@136417.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@136417.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@136417.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@136417.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@136417.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@136431.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@136431.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@136431.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@136431.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@136431.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@136431.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@136445.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@136445.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@136445.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@136445.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@136445.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@136445.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@136459.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@136459.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@136459.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@136459.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@136459.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@136459.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@136473.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@136473.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@136473.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@136473.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@136473.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@136473.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@136487.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@136487.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@136487.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@136487.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@136487.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@136487.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@136501.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@136501.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@136501.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@136501.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@136501.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@136501.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@136515.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@136515.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@136515.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@136515.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@136515.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@136515.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@136529.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@136529.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@136529.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@136529.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@136529.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@136529.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@136543.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@136543.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@136543.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@136543.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@136543.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@136543.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@136557.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@136557.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@136557.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@136557.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@136557.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@136557.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@136571.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@136571.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@136571.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@136571.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@136571.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@136571.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@136585.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@136585.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@136585.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@136585.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@136585.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@136585.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@136599.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@136599.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@136599.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@136599.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@136599.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@136599.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@136613.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@136613.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@136613.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@136613.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@136613.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@136613.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@136627.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@136627.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@136627.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@136627.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@136627.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@136627.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@136641.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@136641.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@136641.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@136641.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@136641.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@136641.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@136655.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@136655.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@136655.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@136655.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@136655.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@136655.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@136669.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@136669.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@136669.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@136669.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@136669.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@136669.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@136683.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@136683.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@136683.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@136683.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@136683.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@136683.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@136697.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@136697.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@136697.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@136697.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@136697.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@136697.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@136711.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@136711.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@136711.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@136711.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@136711.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@136711.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@136725.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@136725.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@136725.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@136725.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@136725.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@136725.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@136739.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@136739.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@136739.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@136739.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@136739.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@136739.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@136753.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@136753.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@136753.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@136753.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@136753.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@136753.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@136767.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@136767.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@136767.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@136767.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@136767.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@136767.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@136781.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@136781.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@136781.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@136781.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@136781.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@136781.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@136795.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@136795.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@136795.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@136795.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@136795.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@136795.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@136809.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@136809.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@136809.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@136809.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@136809.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@136809.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@136823.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@136823.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@136823.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@136823.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@136823.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@136823.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@136837.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@136837.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@136837.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@136837.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@136837.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@136837.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@136851.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@136851.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@136851.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@136851.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@136851.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@136851.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@136865.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@136865.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@136865.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@136865.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@136865.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@136865.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@136879.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@136879.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@136879.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@136879.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@136879.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@136879.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@136893.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@136893.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@136893.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@136893.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@136893.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@136893.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@136907.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@136907.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@136907.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@136907.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@136907.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@136907.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@136921.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@136921.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@136921.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@136921.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@136921.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@136921.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@136935.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@136935.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@136935.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@136935.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@136935.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@136935.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@136949.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@136949.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@136949.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@136949.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@136949.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@136949.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@136963.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@136963.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@136963.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@136963.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@136963.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@136963.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@136977.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@136977.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@136977.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@136977.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@136977.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@136977.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@136991.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@136991.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@136991.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@136991.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@136991.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@136991.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@137005.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@137005.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@137005.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@137005.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@137005.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@137005.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@137019.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@137019.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@137019.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@137019.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@137019.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@137019.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@137033.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@137033.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@137033.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@137033.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@137033.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@137033.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@137047.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@137047.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@137047.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@137047.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@137047.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@137047.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@137061.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@137061.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@137061.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@137061.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@137061.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@137061.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@137075.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@137075.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@137075.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@137075.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@137075.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@137075.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@137089.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@137089.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@137089.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@137089.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@137089.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@137089.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@137103.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@137103.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@137103.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@137103.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@137103.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@137103.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@137117.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@137117.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@137117.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@137117.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@137117.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@137117.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@137131.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@137131.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@137131.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@137131.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@137131.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@137131.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@137145.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@137145.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@137145.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@137145.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@137145.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@137145.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@137159.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@137159.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@137159.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@137159.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@137159.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@137159.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@137173.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@137173.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@137173.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@137173.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@137173.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@137173.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@137187.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@137187.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@137187.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@137187.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@137187.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@137187.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@137201.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@137201.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@137201.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@137201.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@137201.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@137201.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@137215.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@137215.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@137215.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@137215.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@137215.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@137215.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@137229.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@137229.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@137229.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@137229.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@137229.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@137229.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@137243.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@137243.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@137243.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@137243.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@137243.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@137243.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@137257.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@137257.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@137257.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@137257.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@137257.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@137257.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@137271.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@137271.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@137271.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@137271.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@137271.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@137271.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@137285.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@137285.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@137285.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@137285.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@137285.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@137285.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@137299.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@137299.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@137299.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@137299.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@137299.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@137299.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@137313.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@137313.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@137313.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@137313.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@137313.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@137313.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@137327.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@137327.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@137327.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@137327.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@137327.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@137327.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@137341.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@137341.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@137341.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@137341.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@137341.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@137341.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@137355.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@137355.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@137355.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@137355.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@137355.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@137355.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@137369.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@137369.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@137369.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@137369.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@137369.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@137369.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@137383.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@137383.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@137383.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@137383.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@137383.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@137383.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@137397.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@137397.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@137397.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@137397.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@137397.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@137397.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@137411.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@137411.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@137411.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@137411.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@137411.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@137411.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@137425.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@137425.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@137425.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@137425.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@137425.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@137425.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@137439.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@137439.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@137439.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@137439.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@137439.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@137439.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@137453.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@137453.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@137453.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@137453.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@137453.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@137453.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@137467.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@137467.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@137467.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@137467.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@137467.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@137467.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@137481.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@137481.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@137481.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@137481.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@137481.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@137481.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@137495.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@137495.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@137495.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@137495.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@137495.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@137495.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@137509.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@137509.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@137509.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@137509.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@137509.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@137509.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@137523.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@137523.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@137523.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@137523.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@137523.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@137523.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@137537.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@137537.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@137537.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@137537.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@137537.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@137537.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@137551.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@137551.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@137551.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@137551.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@137551.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@137551.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@137565.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@137565.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@137565.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@137565.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@137565.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@137565.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@137579.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@137579.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@137579.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@137579.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@137579.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@137579.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@137593.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@137593.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@137593.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@137593.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@137593.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@137593.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@137607.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@137607.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@137607.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@137607.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@137607.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@137607.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@137621.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@137621.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@137621.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@137621.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@137621.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@137621.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@137635.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@137635.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@137635.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@137635.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@137635.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@137635.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@137649.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@137649.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@137649.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@137649.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@137649.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@137649.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@137663.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@137663.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@137663.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@137663.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@137663.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@137663.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@137677.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@137677.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@137677.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@137677.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@137677.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@137677.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@137691.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@137691.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@137691.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@137691.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@137691.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@137691.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@137705.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@137705.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@137705.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@137705.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@137705.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@137705.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@137719.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@137719.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@137719.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@137719.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@137719.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@137719.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@137733.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@137733.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@137733.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@137733.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@137733.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@137733.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@137747.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@137747.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@137747.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@137747.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@137747.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@137747.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@137761.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@137761.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@137761.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@137761.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@137761.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@137761.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@137775.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@137775.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@137775.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@137775.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@137775.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@137775.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@137789.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@137789.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@137789.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@137789.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@137789.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@137789.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@137803.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@137803.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@137803.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@137803.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@137803.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@137803.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@137817.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@137817.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@137817.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@137817.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@137817.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@137817.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@137831.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@137831.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@137831.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@137831.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@137831.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@137831.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@137845.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@137845.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@137845.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@137845.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@137845.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@137845.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@137859.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@137859.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@137859.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@137859.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@137859.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@137859.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@137873.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@137873.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@137873.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@137873.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@137873.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@137873.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@137887.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@137887.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@137887.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@137887.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@137887.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@137887.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@137901.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@137901.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@137901.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@137901.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@137901.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@137901.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@137915.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@137915.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@137915.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@137915.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@137915.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@137915.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@137929.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@137929.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@137929.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@137929.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@137929.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@137929.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@137943.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@137943.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@137943.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@137943.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@137943.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@137943.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@137957.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@137957.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@137957.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@137957.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@137957.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@137957.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@137971.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@137971.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@137971.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@137971.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@137971.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@137971.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@137985.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@137985.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@137985.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@137985.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@137985.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@137985.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@137999.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@137999.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@137999.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@137999.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@137999.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@137999.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@138013.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@138013.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@138013.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@138013.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@138013.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@138013.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@138027.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@138027.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@138027.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@138027.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@138027.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@138027.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@138041.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@138041.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@138041.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@138041.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@138041.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@138041.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@138055.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@138055.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@138055.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@138055.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@138055.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@138055.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@138069.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@138069.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@138069.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@138069.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@138069.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@138069.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@138083.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@138083.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@138083.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@138083.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@138083.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@138083.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@138097.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@138097.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@138097.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@138097.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@138097.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@138097.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@138111.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@138111.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@138111.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@138111.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@138111.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@138111.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@138125.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@138125.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@138125.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@138125.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@138125.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@138125.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@138139.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@138139.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@138139.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@138139.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@138139.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@138139.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@138153.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@138153.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@138153.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@138153.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@138153.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@138153.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@138167.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@138167.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@138167.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@138167.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@138167.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@138167.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@138181.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@138181.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@138181.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@138181.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@138181.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@138181.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@138195.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@138195.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@138195.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@138195.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@138195.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@138195.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@138209.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@138209.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@138209.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@138209.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@138209.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@138209.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@138223.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@138223.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@138223.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@138223.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@138223.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@138223.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@138237.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@138237.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@138237.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@138237.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@138237.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@138237.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@138251.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@138251.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@138251.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@138251.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@138251.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@138251.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@138265.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@138265.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@138265.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@138265.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@138265.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@138265.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@138279.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@138279.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@138279.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@138279.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@138279.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@138279.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@138293.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@138293.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@138293.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@138293.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@138293.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@138293.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@138307.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@138307.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@138307.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@138307.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@138307.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@138307.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@138321.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@138321.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@138321.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@138321.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@138321.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@138321.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@138335.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@138335.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@138335.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@138335.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@138335.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@138335.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@138349.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@138349.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@138349.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@138349.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@138349.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@138349.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@138363.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@138363.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@138363.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@138363.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@138363.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@138363.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@138377.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@138377.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@138377.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@138377.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@138377.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@138377.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@138391.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@138391.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@138391.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@138391.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@138391.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@138391.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@138405.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@138405.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@138405.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@138405.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@138405.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@138405.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@138419.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@138419.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@138419.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@138419.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@138419.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@138419.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@138433.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@138433.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@138433.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@138433.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@138433.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@138433.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@138447.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@138447.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@138447.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@138447.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@138447.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@138447.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@138461.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@138461.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@138461.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@138461.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@138461.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@138461.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@138475.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@138475.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@138475.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@138475.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@138475.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@138475.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@138489.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@138489.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@138489.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@138489.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@138489.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@138489.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@138503.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@138503.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@138503.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@138503.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@138503.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@138503.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@138517.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@138517.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@138517.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@138517.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@138517.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@138517.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@138531.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@138531.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@138531.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@138531.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@138531.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@138531.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@138545.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@138545.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@138545.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@138545.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@138545.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@138545.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@138559.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@138559.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@138559.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@138559.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@138559.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@138559.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@138573.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@138573.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@138573.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@138573.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@138573.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@138573.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@138587.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@138587.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@138587.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@138587.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@138587.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@138587.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@138601.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@138601.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@138601.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@138601.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@138601.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@138601.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@138615.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@138615.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@138615.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@138615.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@138615.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@138615.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@138629.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@138629.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@138629.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@138629.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@138629.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@138629.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@138643.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@138643.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@138643.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@138643.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@138643.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@138643.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@138657.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@138657.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@138657.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@138657.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@138657.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@138657.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@138671.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@138671.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@138671.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@138671.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@138671.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@138671.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@138685.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@138685.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@138685.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@138685.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@138685.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@138685.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@138699.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@138699.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@138699.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@138699.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@138699.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@138699.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@138713.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@138713.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@138713.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@138713.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@138713.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@138713.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@138727.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@138727.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@138727.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@138727.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@138727.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@138727.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@138741.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@138741.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@138741.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@138741.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@138741.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@138741.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@138755.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@138755.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@138755.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@138755.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@138755.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@138755.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@138769.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@138769.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@138769.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@138769.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@138769.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@138769.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@138783.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@138783.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@138783.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@138783.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@138783.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@138783.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@138797.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@138797.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@138797.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@138797.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@138797.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@138797.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@138811.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@138811.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@138811.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@138811.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@138811.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@138811.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@138825.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@138825.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@138825.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@138825.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@138825.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@138825.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@138839.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@138839.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@138839.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@138839.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@138839.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@138839.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@138853.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@138853.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@138853.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@138853.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@138853.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@138853.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@138867.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@138867.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@138867.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@138867.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@138867.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@138867.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@138881.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@138881.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@138881.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@138881.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@138881.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@138881.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@138895.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@138895.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@138895.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@138895.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@138895.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@138895.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@138909.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@138909.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@138909.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@138909.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@138909.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@138909.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@138923.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@138923.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@138923.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@138923.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@138923.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@138923.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@138937.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@138937.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@138937.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@138937.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@138937.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@138937.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@138951.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@138951.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@138951.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@138951.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@138951.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@138951.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@138965.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@138965.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@138965.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@138965.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@138965.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@138965.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@138979.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@138979.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@138979.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@138979.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@138979.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@138979.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@138993.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@138993.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@138993.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@138993.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@138993.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@138993.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@139007.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@139007.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@139007.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@139007.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@139007.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@139007.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@139021.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@139021.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@139021.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@139021.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@139021.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@139021.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@139035.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@139035.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@139035.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@139035.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@139035.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@139035.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@139049.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@139049.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@139049.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@139049.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@139049.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@139049.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@139063.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@139063.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@139063.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@139063.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@139063.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@139063.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@139077.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@139077.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@139077.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@139077.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@139077.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@139077.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@139091.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@139091.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@139091.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@139091.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@139091.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@139091.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@139105.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@139105.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@139105.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@139105.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@139105.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@139105.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@139119.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@139119.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@139119.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@139119.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@139119.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@139119.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@139133.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@139133.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@139133.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@139133.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@139133.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@139133.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@139147.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@139147.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@139147.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@139147.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@139147.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@139147.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@139161.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@139161.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@139161.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@139161.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@139161.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@139161.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@139175.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@139175.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@139175.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@139175.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@139175.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@139175.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@139189.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@139189.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@139189.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@139189.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@139189.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@139189.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@139203.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@139203.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@139203.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@139203.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@139203.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@139203.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@139217.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@139217.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@139217.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@139217.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@139217.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@139217.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@139231.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@139231.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@139231.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@139231.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@139231.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@139231.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@139245.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@139245.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@139245.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@139245.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@139245.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@139245.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@139259.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@139259.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@139259.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@139259.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@139259.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@139259.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@139273.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@139273.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@139273.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@139273.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@139273.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@139273.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@139287.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@139287.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@139287.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@139287.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@139287.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@139287.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@139301.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@139301.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@139301.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@139301.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@139301.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@139301.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@139315.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@139315.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@139315.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@139315.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@139315.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@139315.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@139329.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@139329.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@139329.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@139329.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@139329.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@139329.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@139343.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@139343.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@139343.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@139343.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@139343.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@139343.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@139357.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@139357.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@139357.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@139357.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@139357.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@139357.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@139371.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@139371.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@139371.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@139371.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@139371.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@139371.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@139385.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@139385.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@139385.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@139385.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@139385.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@139385.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@139399.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@139399.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@139399.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@139399.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@139399.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@139399.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@139413.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@139413.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@139413.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@139413.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@139413.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@139413.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@139427.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@139427.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@139427.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@139427.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@139427.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@139427.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@139441.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@139441.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@139441.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@139441.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@139441.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@139441.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@139455.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@139455.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@139455.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@139455.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@139455.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@139455.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@139469.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@139469.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@139469.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@139469.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@139469.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@139469.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@139483.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@139483.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@139483.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@139483.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@139483.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@139483.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@139497.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@139497.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@139497.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@139497.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@139497.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@139497.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@139511.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@139511.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@139511.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@139511.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@139511.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@139511.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@139525.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@139525.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@139525.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@139525.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@139525.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@139525.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@139539.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@139539.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@139539.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@139539.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@139539.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@139539.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@139553.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@139553.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@139553.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@139553.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@139553.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@139553.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@139567.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@139567.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@139567.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@139567.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@139567.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@139567.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@139581.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@139581.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@139581.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@139581.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@139581.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@139581.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@139595.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@139595.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@139595.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@139595.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@139595.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@139595.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@139609.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@139609.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@139609.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@139609.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@139609.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@139609.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@139623.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@139623.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@139623.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@139623.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@139623.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@139623.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@139637.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@139637.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@139637.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@139637.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@139637.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@139637.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@139651.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@139651.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@139651.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@139651.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@139651.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@139651.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@139665.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@139665.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@139665.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@139665.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@139665.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@139665.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@139679.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@139679.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@139679.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@139679.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@139679.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@139679.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@139693.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@139693.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@139693.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@139693.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@139693.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@139693.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@139707.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@139707.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@139707.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@139707.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@139707.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@139707.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@139721.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@139721.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@139721.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@139721.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@139721.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@139721.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@139735.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@139735.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@139735.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@139735.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@139735.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@139735.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@139749.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@139749.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@139749.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@139749.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@139749.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@139749.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@139763.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@139763.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@139763.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@139763.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@139763.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@139763.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@139777.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@139777.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@139777.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@139777.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@139777.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@139777.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@139791.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@139791.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@139791.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@139791.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@139791.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@139791.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@139805.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@139805.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@139805.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@139805.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@139805.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@139805.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@139819.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@139819.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@139819.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@139819.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@139819.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@139819.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@139833.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@139833.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@139833.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@139833.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@139833.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@139833.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@139847.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@139847.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@139847.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@139847.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@139847.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@139847.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@139861.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@139861.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@139861.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@139861.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@139861.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@139861.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@139875.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@139875.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@139875.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@139875.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@139875.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@139875.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@139889.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@139889.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@139889.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@139889.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@139889.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@139889.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@139903.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@139903.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@139903.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@139903.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@139903.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@139903.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@139917.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@139917.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@139917.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@139917.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@139917.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@139917.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@139931.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@139931.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@139931.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@139931.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@139931.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@139931.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@139945.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@139945.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@139945.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@139945.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@139945.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@139945.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@139959.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@139959.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@139959.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@139959.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@139959.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@139959.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@139973.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@139973.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@139973.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@139973.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@139973.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@139973.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@139987.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@139987.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@139987.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@139987.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@139987.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@139987.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@140001.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@140001.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@140001.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@140001.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@140001.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@140001.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@140015.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@140015.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@140015.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@140015.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@140015.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@140015.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@140029.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@140029.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@140029.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@140029.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@140029.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@140029.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@140043.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@140043.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@140043.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@140043.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@140043.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@140043.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@140057.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@140057.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@140057.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@140057.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@140057.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@140057.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@140071.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@140071.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@140071.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@140071.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@140071.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@140071.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@140085.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@140085.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@140085.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@140085.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@140085.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@140085.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@140099.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@140099.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@140099.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@140099.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@140099.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@140099.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@140113.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@140113.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@140113.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@140113.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@140113.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@140113.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@140127.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@140127.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@140127.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@140127.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@140127.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@140127.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@140141.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@140141.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@140141.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@140141.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@140141.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@140141.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@140155.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@140155.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@140155.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@140155.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@140155.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@140155.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@140169.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@140169.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@140169.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@140169.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@140169.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@140169.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@140183.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@140183.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@140183.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@140183.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@140183.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@140183.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@140197.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@140197.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@140197.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@140197.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@140197.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@140197.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@140211.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@140211.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@140211.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@140211.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@140211.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@140211.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@140225.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@140225.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@140225.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@140225.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@140225.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@140225.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@140239.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@140239.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@140239.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@140239.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@140239.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@140239.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@140253.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@140253.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@140253.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@140253.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@140253.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@140253.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@140267.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@140267.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@140267.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@140267.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@140267.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@140267.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@140281.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@140281.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@140281.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@140281.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@140281.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@140281.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@140295.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@140295.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@140295.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@140295.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@140295.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@140295.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@140309.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@140309.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@140309.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@140309.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@140309.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@140309.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@140323.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@140323.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@140323.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@140323.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@140323.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@140323.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@140337.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@140337.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@140337.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@140337.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@140337.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@140337.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@140351.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@140351.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@140351.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@140351.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@140351.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@140351.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@140365.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@140365.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@140365.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@140365.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@140365.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@140365.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@140379.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@140379.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@140379.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@140379.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@140379.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@140379.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@140393.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@140393.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@140393.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@140393.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@140393.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@140393.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@140407.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@140407.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@140407.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@140407.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@140407.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@140407.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@140421.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@140421.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@140421.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@140421.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@140421.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@140421.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@140435.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@140435.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@140435.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@140435.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@140435.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@140435.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@140449.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@140449.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@140449.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@140449.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@140449.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@140449.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@140463.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@140463.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@140463.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@140463.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@140463.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@140463.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@140477.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@140477.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@140477.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@140477.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@140477.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@140477.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@140491.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@140491.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@140491.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@140491.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@140491.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@140491.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@140505.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@140505.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@140505.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@140505.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@140505.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@140505.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@140519.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@140519.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@140519.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@140519.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@140519.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@140519.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@140533.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@140533.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@140533.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@140533.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@140533.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@140533.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@140547.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@140547.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@140547.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@140547.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@140547.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@140547.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@140561.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@140561.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@140561.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@140561.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@140561.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@140561.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@140575.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@140575.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@140575.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@140575.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@140575.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@140575.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@140589.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@140589.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@140589.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@140589.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@140589.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@140589.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@140603.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@140603.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@140603.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@140603.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@140603.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@140603.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@140617.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@140617.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@140617.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@140617.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@140617.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@140617.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@140631.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@140631.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@140631.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@140631.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@140631.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@140631.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@140645.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@140645.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@140645.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@140645.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@140645.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@140645.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@140659.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@140659.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@140659.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@140659.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@140659.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@140659.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@140673.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@140673.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@140673.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@140673.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@140673.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@140673.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@140687.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@140687.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@140687.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@133649.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@133661.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@133662.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@133680.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@133692.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@133704.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@133705.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@133646.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@133658.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@133677.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@133689.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@133701.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@133715.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@133729.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@133743.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@133757.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@133771.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@133785.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@133799.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@133813.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@133827.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@133841.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@133855.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@133869.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@133883.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@133897.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@133911.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@133925.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@133939.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@133953.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@133967.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@133981.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@133995.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@134009.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@134023.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@134037.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@134051.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@134065.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@134079.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@134093.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@134107.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@134121.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@134135.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@134149.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@134163.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@134177.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@134191.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@134205.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@134219.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@134233.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@134247.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@134261.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@134275.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@134289.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@134303.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@134317.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@134331.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@134345.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@134359.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@134373.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@134387.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@134401.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@134415.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@134429.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@134443.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@134457.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@134471.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@134485.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@134499.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@134513.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@134527.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@134541.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@134555.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@134569.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@134583.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@134597.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@134611.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@134625.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@134639.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@134653.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@134667.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@134681.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@134695.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@134709.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@134723.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@134737.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@134751.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@134765.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@134779.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@134793.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@134807.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@134821.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@134835.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@134849.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@134863.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@134877.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@134891.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@134905.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@134919.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@134933.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@134947.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@134961.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@134975.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@134989.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@135003.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@135017.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@135031.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@135045.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@135059.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@135073.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@135087.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@135101.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@135115.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@135129.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@135143.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@135157.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@135171.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@135185.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@135199.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@135213.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@135227.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@135241.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@135255.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@135269.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@135283.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@135297.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@135311.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@135325.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@135339.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@135353.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@135367.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@135381.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@135395.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@135409.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@135423.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@135437.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@135451.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@135465.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@135479.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@135493.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@135507.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@135521.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@135535.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@135549.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@135563.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@135577.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@135591.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@135605.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@135619.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@135633.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@135647.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@135661.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@135675.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@135689.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@135703.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@135717.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@135731.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@135745.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@135759.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@135773.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@135787.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@135801.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@135815.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@135829.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@135843.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@135857.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@135871.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@135885.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@135899.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@135913.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@135927.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@135941.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@135955.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@135969.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@135983.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@135997.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@136011.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@136025.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@136039.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@136053.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@136067.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@136081.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@136095.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@136109.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@136123.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@136137.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@136151.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@136165.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@136179.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@136193.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@136207.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@136221.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@136235.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@136249.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@136263.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@136277.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@136291.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@136305.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@136319.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@136333.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@136347.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@136361.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@136375.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@136389.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@136403.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@136417.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@136431.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@136445.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@136459.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@136473.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@136487.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@136501.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@136515.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@136529.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@136543.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@136557.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@136571.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@136585.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@136599.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@136613.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@136627.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@136641.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@136655.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@136669.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@136683.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@136697.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@136711.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@136725.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@136739.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@136753.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@136767.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@136781.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@136795.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@136809.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@136823.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@136837.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@136851.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@136865.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@136879.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@136893.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@136907.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@136921.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@136935.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@136949.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@136963.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@136977.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@136991.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@137005.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@137019.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@137033.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@137047.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@137061.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@137075.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@137089.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@137103.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@137117.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@137131.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@137145.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@137159.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@137173.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@137187.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@137201.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@137215.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@137229.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@137243.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@137257.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@137271.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@137285.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@137299.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@137313.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@137327.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@137341.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@137355.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@137369.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@137383.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@137397.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@137411.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@137425.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@137439.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@137453.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@137467.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@137481.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@137495.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@137509.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@137523.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@137537.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@137551.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@137565.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@137579.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@137593.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@137607.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@137621.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@137635.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@137649.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@137663.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@137677.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@137691.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@137705.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@137719.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@137733.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@137747.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@137761.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@137775.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@137789.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@137803.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@137817.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@137831.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@137845.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@137859.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@137873.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@137887.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@137901.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@137915.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@137929.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@137943.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@137957.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@137971.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@137985.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@137999.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@138013.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@138027.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@138041.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@138055.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@138069.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@138083.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@138097.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@138111.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@138125.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@138139.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@138153.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@138167.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@138181.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@138195.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@138209.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@138223.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@138237.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@138251.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@138265.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@138279.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@138293.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@138307.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@138321.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@138335.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@138349.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@138363.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@138377.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@138391.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@138405.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@138419.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@138433.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@138447.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@138461.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@138475.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@138489.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@138503.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@138517.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@138531.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@138545.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@138559.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@138573.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@138587.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@138601.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@138615.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@138629.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@138643.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@138657.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@138671.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@138685.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@138699.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@138713.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@138727.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@138741.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@138755.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@138769.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@138783.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@138797.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@138811.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@138825.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@138839.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@138853.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@138867.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@138881.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@138895.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@138909.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@138923.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@138937.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@138951.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@138965.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@138979.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@138993.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@139007.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@139021.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@139035.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@139049.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@139063.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@139077.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@139091.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@139105.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@139119.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@139133.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@139147.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@139161.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@139175.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@139189.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@139203.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@139217.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@139231.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@139245.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@139259.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@139273.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@139287.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@139301.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@139315.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@139329.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@139343.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@139357.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@139371.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@139385.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@139399.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@139413.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@139427.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@139441.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@139455.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@139469.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@139483.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@139497.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@139511.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@139525.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@139539.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@139553.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@139567.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@139581.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@139595.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@139609.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@139623.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@139637.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@139651.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@139665.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@139679.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@139693.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@139707.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@139721.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@139735.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@139749.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@139763.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@139777.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@139791.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@139805.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@139819.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@139833.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@139847.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@139861.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@139875.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@139889.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@139903.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@139917.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@139931.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@139945.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@139959.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@139973.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@139987.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@140001.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@140015.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@140029.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@140043.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@140057.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@140071.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@140085.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@140099.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@140113.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@140127.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@140141.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@140155.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@140169.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@140183.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@140197.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@140211.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@140225.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@140239.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@140253.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@140267.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@140281.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@140295.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@140309.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@140323.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@140337.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@140351.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@140365.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@140379.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@140393.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@140407.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@140421.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@140435.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@140449.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@140463.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@140477.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@140491.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@140505.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@140519.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@140533.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@140547.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@140561.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@140575.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@140589.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@140603.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@140617.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@140631.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@140645.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@140659.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@140673.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@140687.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@133649.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@133661.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@133662.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@133680.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@133692.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@133704.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@133705.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@141698.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@141704.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@141705.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@141706.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@141707.4]
  assign regs_0_clock = clock; // @[:@133647.4]
  assign regs_0_reset = reset; // @[:@133648.4 RegFile.scala 82:16:@133654.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@133652.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@133656.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@133651.4]
  assign regs_1_clock = clock; // @[:@133659.4]
  assign regs_1_reset = reset; // @[:@133660.4 RegFile.scala 70:16:@133672.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@133670.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@133675.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@133666.4]
  assign regs_2_clock = clock; // @[:@133678.4]
  assign regs_2_reset = reset; // @[:@133679.4 RegFile.scala 82:16:@133685.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@133683.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@133687.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@133682.4]
  assign regs_3_clock = clock; // @[:@133690.4]
  assign regs_3_reset = reset; // @[:@133691.4 RegFile.scala 82:16:@133697.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@133695.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@133699.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@133694.4]
  assign regs_4_clock = clock; // @[:@133702.4]
  assign regs_4_reset = io_reset; // @[:@133703.4 RegFile.scala 76:16:@133710.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@133709.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@133713.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@133707.4]
  assign regs_5_clock = clock; // @[:@133716.4]
  assign regs_5_reset = io_reset; // @[:@133717.4 RegFile.scala 76:16:@133724.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@133723.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@133727.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@133721.4]
  assign regs_6_clock = clock; // @[:@133730.4]
  assign regs_6_reset = io_reset; // @[:@133731.4 RegFile.scala 76:16:@133738.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@133737.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@133741.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@133735.4]
  assign regs_7_clock = clock; // @[:@133744.4]
  assign regs_7_reset = io_reset; // @[:@133745.4 RegFile.scala 76:16:@133752.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@133751.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@133755.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@133749.4]
  assign regs_8_clock = clock; // @[:@133758.4]
  assign regs_8_reset = io_reset; // @[:@133759.4 RegFile.scala 76:16:@133766.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@133765.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@133769.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@133763.4]
  assign regs_9_clock = clock; // @[:@133772.4]
  assign regs_9_reset = io_reset; // @[:@133773.4 RegFile.scala 76:16:@133780.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@133779.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@133783.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@133777.4]
  assign regs_10_clock = clock; // @[:@133786.4]
  assign regs_10_reset = io_reset; // @[:@133787.4 RegFile.scala 76:16:@133794.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@133793.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@133797.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@133791.4]
  assign regs_11_clock = clock; // @[:@133800.4]
  assign regs_11_reset = io_reset; // @[:@133801.4 RegFile.scala 76:16:@133808.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@133807.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@133811.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@133805.4]
  assign regs_12_clock = clock; // @[:@133814.4]
  assign regs_12_reset = io_reset; // @[:@133815.4 RegFile.scala 76:16:@133822.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@133821.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@133825.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@133819.4]
  assign regs_13_clock = clock; // @[:@133828.4]
  assign regs_13_reset = io_reset; // @[:@133829.4 RegFile.scala 76:16:@133836.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@133835.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@133839.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@133833.4]
  assign regs_14_clock = clock; // @[:@133842.4]
  assign regs_14_reset = io_reset; // @[:@133843.4 RegFile.scala 76:16:@133850.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@133849.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@133853.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@133847.4]
  assign regs_15_clock = clock; // @[:@133856.4]
  assign regs_15_reset = io_reset; // @[:@133857.4 RegFile.scala 76:16:@133864.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@133863.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@133867.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@133861.4]
  assign regs_16_clock = clock; // @[:@133870.4]
  assign regs_16_reset = io_reset; // @[:@133871.4 RegFile.scala 76:16:@133878.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@133877.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@133881.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@133875.4]
  assign regs_17_clock = clock; // @[:@133884.4]
  assign regs_17_reset = io_reset; // @[:@133885.4 RegFile.scala 76:16:@133892.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@133891.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@133895.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@133889.4]
  assign regs_18_clock = clock; // @[:@133898.4]
  assign regs_18_reset = io_reset; // @[:@133899.4 RegFile.scala 76:16:@133906.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@133905.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@133909.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@133903.4]
  assign regs_19_clock = clock; // @[:@133912.4]
  assign regs_19_reset = io_reset; // @[:@133913.4 RegFile.scala 76:16:@133920.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@133919.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@133923.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@133917.4]
  assign regs_20_clock = clock; // @[:@133926.4]
  assign regs_20_reset = io_reset; // @[:@133927.4 RegFile.scala 76:16:@133934.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@133933.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@133937.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@133931.4]
  assign regs_21_clock = clock; // @[:@133940.4]
  assign regs_21_reset = io_reset; // @[:@133941.4 RegFile.scala 76:16:@133948.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@133947.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@133951.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@133945.4]
  assign regs_22_clock = clock; // @[:@133954.4]
  assign regs_22_reset = io_reset; // @[:@133955.4 RegFile.scala 76:16:@133962.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@133961.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@133965.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@133959.4]
  assign regs_23_clock = clock; // @[:@133968.4]
  assign regs_23_reset = io_reset; // @[:@133969.4 RegFile.scala 76:16:@133976.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@133975.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@133979.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@133973.4]
  assign regs_24_clock = clock; // @[:@133982.4]
  assign regs_24_reset = io_reset; // @[:@133983.4 RegFile.scala 76:16:@133990.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@133989.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@133993.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@133987.4]
  assign regs_25_clock = clock; // @[:@133996.4]
  assign regs_25_reset = io_reset; // @[:@133997.4 RegFile.scala 76:16:@134004.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@134003.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@134007.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@134001.4]
  assign regs_26_clock = clock; // @[:@134010.4]
  assign regs_26_reset = io_reset; // @[:@134011.4 RegFile.scala 76:16:@134018.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@134017.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@134021.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@134015.4]
  assign regs_27_clock = clock; // @[:@134024.4]
  assign regs_27_reset = io_reset; // @[:@134025.4 RegFile.scala 76:16:@134032.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@134031.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@134035.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@134029.4]
  assign regs_28_clock = clock; // @[:@134038.4]
  assign regs_28_reset = io_reset; // @[:@134039.4 RegFile.scala 76:16:@134046.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@134045.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@134049.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@134043.4]
  assign regs_29_clock = clock; // @[:@134052.4]
  assign regs_29_reset = io_reset; // @[:@134053.4 RegFile.scala 76:16:@134060.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@134059.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@134063.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@134057.4]
  assign regs_30_clock = clock; // @[:@134066.4]
  assign regs_30_reset = io_reset; // @[:@134067.4 RegFile.scala 76:16:@134074.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@134073.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@134077.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@134071.4]
  assign regs_31_clock = clock; // @[:@134080.4]
  assign regs_31_reset = io_reset; // @[:@134081.4 RegFile.scala 76:16:@134088.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@134087.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@134091.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@134085.4]
  assign regs_32_clock = clock; // @[:@134094.4]
  assign regs_32_reset = io_reset; // @[:@134095.4 RegFile.scala 76:16:@134102.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@134101.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@134105.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@134099.4]
  assign regs_33_clock = clock; // @[:@134108.4]
  assign regs_33_reset = io_reset; // @[:@134109.4 RegFile.scala 76:16:@134116.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@134115.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@134119.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@134113.4]
  assign regs_34_clock = clock; // @[:@134122.4]
  assign regs_34_reset = io_reset; // @[:@134123.4 RegFile.scala 76:16:@134130.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@134129.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@134133.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@134127.4]
  assign regs_35_clock = clock; // @[:@134136.4]
  assign regs_35_reset = io_reset; // @[:@134137.4 RegFile.scala 76:16:@134144.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@134143.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@134147.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@134141.4]
  assign regs_36_clock = clock; // @[:@134150.4]
  assign regs_36_reset = io_reset; // @[:@134151.4 RegFile.scala 76:16:@134158.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@134157.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@134161.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@134155.4]
  assign regs_37_clock = clock; // @[:@134164.4]
  assign regs_37_reset = io_reset; // @[:@134165.4 RegFile.scala 76:16:@134172.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@134171.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@134175.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@134169.4]
  assign regs_38_clock = clock; // @[:@134178.4]
  assign regs_38_reset = io_reset; // @[:@134179.4 RegFile.scala 76:16:@134186.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@134185.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@134189.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@134183.4]
  assign regs_39_clock = clock; // @[:@134192.4]
  assign regs_39_reset = io_reset; // @[:@134193.4 RegFile.scala 76:16:@134200.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@134199.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@134203.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@134197.4]
  assign regs_40_clock = clock; // @[:@134206.4]
  assign regs_40_reset = io_reset; // @[:@134207.4 RegFile.scala 76:16:@134214.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@134213.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@134217.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@134211.4]
  assign regs_41_clock = clock; // @[:@134220.4]
  assign regs_41_reset = io_reset; // @[:@134221.4 RegFile.scala 76:16:@134228.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@134227.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@134231.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@134225.4]
  assign regs_42_clock = clock; // @[:@134234.4]
  assign regs_42_reset = io_reset; // @[:@134235.4 RegFile.scala 76:16:@134242.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@134241.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@134245.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@134239.4]
  assign regs_43_clock = clock; // @[:@134248.4]
  assign regs_43_reset = io_reset; // @[:@134249.4 RegFile.scala 76:16:@134256.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@134255.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@134259.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@134253.4]
  assign regs_44_clock = clock; // @[:@134262.4]
  assign regs_44_reset = io_reset; // @[:@134263.4 RegFile.scala 76:16:@134270.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@134269.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@134273.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@134267.4]
  assign regs_45_clock = clock; // @[:@134276.4]
  assign regs_45_reset = io_reset; // @[:@134277.4 RegFile.scala 76:16:@134284.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@134283.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@134287.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@134281.4]
  assign regs_46_clock = clock; // @[:@134290.4]
  assign regs_46_reset = io_reset; // @[:@134291.4 RegFile.scala 76:16:@134298.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@134297.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@134301.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@134295.4]
  assign regs_47_clock = clock; // @[:@134304.4]
  assign regs_47_reset = io_reset; // @[:@134305.4 RegFile.scala 76:16:@134312.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@134311.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@134315.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@134309.4]
  assign regs_48_clock = clock; // @[:@134318.4]
  assign regs_48_reset = io_reset; // @[:@134319.4 RegFile.scala 76:16:@134326.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@134325.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@134329.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@134323.4]
  assign regs_49_clock = clock; // @[:@134332.4]
  assign regs_49_reset = io_reset; // @[:@134333.4 RegFile.scala 76:16:@134340.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@134339.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@134343.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@134337.4]
  assign regs_50_clock = clock; // @[:@134346.4]
  assign regs_50_reset = io_reset; // @[:@134347.4 RegFile.scala 76:16:@134354.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@134353.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@134357.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@134351.4]
  assign regs_51_clock = clock; // @[:@134360.4]
  assign regs_51_reset = io_reset; // @[:@134361.4 RegFile.scala 76:16:@134368.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@134367.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@134371.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@134365.4]
  assign regs_52_clock = clock; // @[:@134374.4]
  assign regs_52_reset = io_reset; // @[:@134375.4 RegFile.scala 76:16:@134382.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@134381.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@134385.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@134379.4]
  assign regs_53_clock = clock; // @[:@134388.4]
  assign regs_53_reset = io_reset; // @[:@134389.4 RegFile.scala 76:16:@134396.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@134395.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@134399.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@134393.4]
  assign regs_54_clock = clock; // @[:@134402.4]
  assign regs_54_reset = io_reset; // @[:@134403.4 RegFile.scala 76:16:@134410.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@134409.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@134413.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@134407.4]
  assign regs_55_clock = clock; // @[:@134416.4]
  assign regs_55_reset = io_reset; // @[:@134417.4 RegFile.scala 76:16:@134424.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@134423.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@134427.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@134421.4]
  assign regs_56_clock = clock; // @[:@134430.4]
  assign regs_56_reset = io_reset; // @[:@134431.4 RegFile.scala 76:16:@134438.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@134437.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@134441.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@134435.4]
  assign regs_57_clock = clock; // @[:@134444.4]
  assign regs_57_reset = io_reset; // @[:@134445.4 RegFile.scala 76:16:@134452.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@134451.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@134455.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@134449.4]
  assign regs_58_clock = clock; // @[:@134458.4]
  assign regs_58_reset = io_reset; // @[:@134459.4 RegFile.scala 76:16:@134466.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@134465.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@134469.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@134463.4]
  assign regs_59_clock = clock; // @[:@134472.4]
  assign regs_59_reset = io_reset; // @[:@134473.4 RegFile.scala 76:16:@134480.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@134479.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@134483.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@134477.4]
  assign regs_60_clock = clock; // @[:@134486.4]
  assign regs_60_reset = io_reset; // @[:@134487.4 RegFile.scala 76:16:@134494.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@134493.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@134497.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@134491.4]
  assign regs_61_clock = clock; // @[:@134500.4]
  assign regs_61_reset = io_reset; // @[:@134501.4 RegFile.scala 76:16:@134508.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@134507.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@134511.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@134505.4]
  assign regs_62_clock = clock; // @[:@134514.4]
  assign regs_62_reset = io_reset; // @[:@134515.4 RegFile.scala 76:16:@134522.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@134521.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@134525.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@134519.4]
  assign regs_63_clock = clock; // @[:@134528.4]
  assign regs_63_reset = io_reset; // @[:@134529.4 RegFile.scala 76:16:@134536.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@134535.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@134539.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@134533.4]
  assign regs_64_clock = clock; // @[:@134542.4]
  assign regs_64_reset = io_reset; // @[:@134543.4 RegFile.scala 76:16:@134550.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@134549.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@134553.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@134547.4]
  assign regs_65_clock = clock; // @[:@134556.4]
  assign regs_65_reset = io_reset; // @[:@134557.4 RegFile.scala 76:16:@134564.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@134563.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@134567.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@134561.4]
  assign regs_66_clock = clock; // @[:@134570.4]
  assign regs_66_reset = io_reset; // @[:@134571.4 RegFile.scala 76:16:@134578.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@134577.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@134581.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@134575.4]
  assign regs_67_clock = clock; // @[:@134584.4]
  assign regs_67_reset = io_reset; // @[:@134585.4 RegFile.scala 76:16:@134592.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@134591.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@134595.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@134589.4]
  assign regs_68_clock = clock; // @[:@134598.4]
  assign regs_68_reset = io_reset; // @[:@134599.4 RegFile.scala 76:16:@134606.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@134605.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@134609.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@134603.4]
  assign regs_69_clock = clock; // @[:@134612.4]
  assign regs_69_reset = io_reset; // @[:@134613.4 RegFile.scala 76:16:@134620.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@134619.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@134623.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@134617.4]
  assign regs_70_clock = clock; // @[:@134626.4]
  assign regs_70_reset = io_reset; // @[:@134627.4 RegFile.scala 76:16:@134634.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@134633.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@134637.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@134631.4]
  assign regs_71_clock = clock; // @[:@134640.4]
  assign regs_71_reset = io_reset; // @[:@134641.4 RegFile.scala 76:16:@134648.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@134647.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@134651.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@134645.4]
  assign regs_72_clock = clock; // @[:@134654.4]
  assign regs_72_reset = io_reset; // @[:@134655.4 RegFile.scala 76:16:@134662.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@134661.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@134665.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@134659.4]
  assign regs_73_clock = clock; // @[:@134668.4]
  assign regs_73_reset = io_reset; // @[:@134669.4 RegFile.scala 76:16:@134676.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@134675.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@134679.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@134673.4]
  assign regs_74_clock = clock; // @[:@134682.4]
  assign regs_74_reset = io_reset; // @[:@134683.4 RegFile.scala 76:16:@134690.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@134689.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@134693.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@134687.4]
  assign regs_75_clock = clock; // @[:@134696.4]
  assign regs_75_reset = io_reset; // @[:@134697.4 RegFile.scala 76:16:@134704.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@134703.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@134707.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@134701.4]
  assign regs_76_clock = clock; // @[:@134710.4]
  assign regs_76_reset = io_reset; // @[:@134711.4 RegFile.scala 76:16:@134718.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@134717.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@134721.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@134715.4]
  assign regs_77_clock = clock; // @[:@134724.4]
  assign regs_77_reset = io_reset; // @[:@134725.4 RegFile.scala 76:16:@134732.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@134731.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@134735.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@134729.4]
  assign regs_78_clock = clock; // @[:@134738.4]
  assign regs_78_reset = io_reset; // @[:@134739.4 RegFile.scala 76:16:@134746.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@134745.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@134749.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@134743.4]
  assign regs_79_clock = clock; // @[:@134752.4]
  assign regs_79_reset = io_reset; // @[:@134753.4 RegFile.scala 76:16:@134760.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@134759.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@134763.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@134757.4]
  assign regs_80_clock = clock; // @[:@134766.4]
  assign regs_80_reset = io_reset; // @[:@134767.4 RegFile.scala 76:16:@134774.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@134773.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@134777.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@134771.4]
  assign regs_81_clock = clock; // @[:@134780.4]
  assign regs_81_reset = io_reset; // @[:@134781.4 RegFile.scala 76:16:@134788.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@134787.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@134791.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@134785.4]
  assign regs_82_clock = clock; // @[:@134794.4]
  assign regs_82_reset = io_reset; // @[:@134795.4 RegFile.scala 76:16:@134802.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@134801.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@134805.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@134799.4]
  assign regs_83_clock = clock; // @[:@134808.4]
  assign regs_83_reset = io_reset; // @[:@134809.4 RegFile.scala 76:16:@134816.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@134815.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@134819.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@134813.4]
  assign regs_84_clock = clock; // @[:@134822.4]
  assign regs_84_reset = io_reset; // @[:@134823.4 RegFile.scala 76:16:@134830.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@134829.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@134833.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@134827.4]
  assign regs_85_clock = clock; // @[:@134836.4]
  assign regs_85_reset = io_reset; // @[:@134837.4 RegFile.scala 76:16:@134844.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@134843.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@134847.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@134841.4]
  assign regs_86_clock = clock; // @[:@134850.4]
  assign regs_86_reset = io_reset; // @[:@134851.4 RegFile.scala 76:16:@134858.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@134857.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@134861.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@134855.4]
  assign regs_87_clock = clock; // @[:@134864.4]
  assign regs_87_reset = io_reset; // @[:@134865.4 RegFile.scala 76:16:@134872.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@134871.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@134875.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@134869.4]
  assign regs_88_clock = clock; // @[:@134878.4]
  assign regs_88_reset = io_reset; // @[:@134879.4 RegFile.scala 76:16:@134886.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@134885.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@134889.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@134883.4]
  assign regs_89_clock = clock; // @[:@134892.4]
  assign regs_89_reset = io_reset; // @[:@134893.4 RegFile.scala 76:16:@134900.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@134899.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@134903.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@134897.4]
  assign regs_90_clock = clock; // @[:@134906.4]
  assign regs_90_reset = io_reset; // @[:@134907.4 RegFile.scala 76:16:@134914.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@134913.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@134917.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@134911.4]
  assign regs_91_clock = clock; // @[:@134920.4]
  assign regs_91_reset = io_reset; // @[:@134921.4 RegFile.scala 76:16:@134928.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@134927.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@134931.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@134925.4]
  assign regs_92_clock = clock; // @[:@134934.4]
  assign regs_92_reset = io_reset; // @[:@134935.4 RegFile.scala 76:16:@134942.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@134941.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@134945.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@134939.4]
  assign regs_93_clock = clock; // @[:@134948.4]
  assign regs_93_reset = io_reset; // @[:@134949.4 RegFile.scala 76:16:@134956.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@134955.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@134959.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@134953.4]
  assign regs_94_clock = clock; // @[:@134962.4]
  assign regs_94_reset = io_reset; // @[:@134963.4 RegFile.scala 76:16:@134970.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@134969.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@134973.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@134967.4]
  assign regs_95_clock = clock; // @[:@134976.4]
  assign regs_95_reset = io_reset; // @[:@134977.4 RegFile.scala 76:16:@134984.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@134983.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@134987.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@134981.4]
  assign regs_96_clock = clock; // @[:@134990.4]
  assign regs_96_reset = io_reset; // @[:@134991.4 RegFile.scala 76:16:@134998.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@134997.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@135001.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@134995.4]
  assign regs_97_clock = clock; // @[:@135004.4]
  assign regs_97_reset = io_reset; // @[:@135005.4 RegFile.scala 76:16:@135012.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@135011.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@135015.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@135009.4]
  assign regs_98_clock = clock; // @[:@135018.4]
  assign regs_98_reset = io_reset; // @[:@135019.4 RegFile.scala 76:16:@135026.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@135025.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@135029.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@135023.4]
  assign regs_99_clock = clock; // @[:@135032.4]
  assign regs_99_reset = io_reset; // @[:@135033.4 RegFile.scala 76:16:@135040.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@135039.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@135043.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@135037.4]
  assign regs_100_clock = clock; // @[:@135046.4]
  assign regs_100_reset = io_reset; // @[:@135047.4 RegFile.scala 76:16:@135054.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@135053.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@135057.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@135051.4]
  assign regs_101_clock = clock; // @[:@135060.4]
  assign regs_101_reset = io_reset; // @[:@135061.4 RegFile.scala 76:16:@135068.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@135067.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@135071.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@135065.4]
  assign regs_102_clock = clock; // @[:@135074.4]
  assign regs_102_reset = io_reset; // @[:@135075.4 RegFile.scala 76:16:@135082.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@135081.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@135085.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@135079.4]
  assign regs_103_clock = clock; // @[:@135088.4]
  assign regs_103_reset = io_reset; // @[:@135089.4 RegFile.scala 76:16:@135096.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@135095.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@135099.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@135093.4]
  assign regs_104_clock = clock; // @[:@135102.4]
  assign regs_104_reset = io_reset; // @[:@135103.4 RegFile.scala 76:16:@135110.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@135109.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@135113.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@135107.4]
  assign regs_105_clock = clock; // @[:@135116.4]
  assign regs_105_reset = io_reset; // @[:@135117.4 RegFile.scala 76:16:@135124.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@135123.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@135127.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@135121.4]
  assign regs_106_clock = clock; // @[:@135130.4]
  assign regs_106_reset = io_reset; // @[:@135131.4 RegFile.scala 76:16:@135138.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@135137.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@135141.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@135135.4]
  assign regs_107_clock = clock; // @[:@135144.4]
  assign regs_107_reset = io_reset; // @[:@135145.4 RegFile.scala 76:16:@135152.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@135151.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@135155.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@135149.4]
  assign regs_108_clock = clock; // @[:@135158.4]
  assign regs_108_reset = io_reset; // @[:@135159.4 RegFile.scala 76:16:@135166.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@135165.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@135169.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@135163.4]
  assign regs_109_clock = clock; // @[:@135172.4]
  assign regs_109_reset = io_reset; // @[:@135173.4 RegFile.scala 76:16:@135180.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@135179.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@135183.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@135177.4]
  assign regs_110_clock = clock; // @[:@135186.4]
  assign regs_110_reset = io_reset; // @[:@135187.4 RegFile.scala 76:16:@135194.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@135193.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@135197.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@135191.4]
  assign regs_111_clock = clock; // @[:@135200.4]
  assign regs_111_reset = io_reset; // @[:@135201.4 RegFile.scala 76:16:@135208.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@135207.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@135211.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@135205.4]
  assign regs_112_clock = clock; // @[:@135214.4]
  assign regs_112_reset = io_reset; // @[:@135215.4 RegFile.scala 76:16:@135222.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@135221.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@135225.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@135219.4]
  assign regs_113_clock = clock; // @[:@135228.4]
  assign regs_113_reset = io_reset; // @[:@135229.4 RegFile.scala 76:16:@135236.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@135235.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@135239.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@135233.4]
  assign regs_114_clock = clock; // @[:@135242.4]
  assign regs_114_reset = io_reset; // @[:@135243.4 RegFile.scala 76:16:@135250.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@135249.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@135253.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@135247.4]
  assign regs_115_clock = clock; // @[:@135256.4]
  assign regs_115_reset = io_reset; // @[:@135257.4 RegFile.scala 76:16:@135264.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@135263.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@135267.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@135261.4]
  assign regs_116_clock = clock; // @[:@135270.4]
  assign regs_116_reset = io_reset; // @[:@135271.4 RegFile.scala 76:16:@135278.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@135277.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@135281.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@135275.4]
  assign regs_117_clock = clock; // @[:@135284.4]
  assign regs_117_reset = io_reset; // @[:@135285.4 RegFile.scala 76:16:@135292.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@135291.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@135295.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@135289.4]
  assign regs_118_clock = clock; // @[:@135298.4]
  assign regs_118_reset = io_reset; // @[:@135299.4 RegFile.scala 76:16:@135306.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@135305.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@135309.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@135303.4]
  assign regs_119_clock = clock; // @[:@135312.4]
  assign regs_119_reset = io_reset; // @[:@135313.4 RegFile.scala 76:16:@135320.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@135319.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@135323.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@135317.4]
  assign regs_120_clock = clock; // @[:@135326.4]
  assign regs_120_reset = io_reset; // @[:@135327.4 RegFile.scala 76:16:@135334.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@135333.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@135337.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@135331.4]
  assign regs_121_clock = clock; // @[:@135340.4]
  assign regs_121_reset = io_reset; // @[:@135341.4 RegFile.scala 76:16:@135348.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@135347.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@135351.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@135345.4]
  assign regs_122_clock = clock; // @[:@135354.4]
  assign regs_122_reset = io_reset; // @[:@135355.4 RegFile.scala 76:16:@135362.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@135361.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@135365.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@135359.4]
  assign regs_123_clock = clock; // @[:@135368.4]
  assign regs_123_reset = io_reset; // @[:@135369.4 RegFile.scala 76:16:@135376.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@135375.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@135379.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@135373.4]
  assign regs_124_clock = clock; // @[:@135382.4]
  assign regs_124_reset = io_reset; // @[:@135383.4 RegFile.scala 76:16:@135390.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@135389.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@135393.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@135387.4]
  assign regs_125_clock = clock; // @[:@135396.4]
  assign regs_125_reset = io_reset; // @[:@135397.4 RegFile.scala 76:16:@135404.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@135403.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@135407.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@135401.4]
  assign regs_126_clock = clock; // @[:@135410.4]
  assign regs_126_reset = io_reset; // @[:@135411.4 RegFile.scala 76:16:@135418.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@135417.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@135421.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@135415.4]
  assign regs_127_clock = clock; // @[:@135424.4]
  assign regs_127_reset = io_reset; // @[:@135425.4 RegFile.scala 76:16:@135432.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@135431.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@135435.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@135429.4]
  assign regs_128_clock = clock; // @[:@135438.4]
  assign regs_128_reset = io_reset; // @[:@135439.4 RegFile.scala 76:16:@135446.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@135445.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@135449.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@135443.4]
  assign regs_129_clock = clock; // @[:@135452.4]
  assign regs_129_reset = io_reset; // @[:@135453.4 RegFile.scala 76:16:@135460.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@135459.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@135463.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@135457.4]
  assign regs_130_clock = clock; // @[:@135466.4]
  assign regs_130_reset = io_reset; // @[:@135467.4 RegFile.scala 76:16:@135474.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@135473.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@135477.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@135471.4]
  assign regs_131_clock = clock; // @[:@135480.4]
  assign regs_131_reset = io_reset; // @[:@135481.4 RegFile.scala 76:16:@135488.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@135487.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@135491.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@135485.4]
  assign regs_132_clock = clock; // @[:@135494.4]
  assign regs_132_reset = io_reset; // @[:@135495.4 RegFile.scala 76:16:@135502.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@135501.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@135505.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@135499.4]
  assign regs_133_clock = clock; // @[:@135508.4]
  assign regs_133_reset = io_reset; // @[:@135509.4 RegFile.scala 76:16:@135516.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@135515.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@135519.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@135513.4]
  assign regs_134_clock = clock; // @[:@135522.4]
  assign regs_134_reset = io_reset; // @[:@135523.4 RegFile.scala 76:16:@135530.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@135529.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@135533.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@135527.4]
  assign regs_135_clock = clock; // @[:@135536.4]
  assign regs_135_reset = io_reset; // @[:@135537.4 RegFile.scala 76:16:@135544.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@135543.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@135547.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@135541.4]
  assign regs_136_clock = clock; // @[:@135550.4]
  assign regs_136_reset = io_reset; // @[:@135551.4 RegFile.scala 76:16:@135558.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@135557.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@135561.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@135555.4]
  assign regs_137_clock = clock; // @[:@135564.4]
  assign regs_137_reset = io_reset; // @[:@135565.4 RegFile.scala 76:16:@135572.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@135571.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@135575.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@135569.4]
  assign regs_138_clock = clock; // @[:@135578.4]
  assign regs_138_reset = io_reset; // @[:@135579.4 RegFile.scala 76:16:@135586.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@135585.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@135589.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@135583.4]
  assign regs_139_clock = clock; // @[:@135592.4]
  assign regs_139_reset = io_reset; // @[:@135593.4 RegFile.scala 76:16:@135600.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@135599.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@135603.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@135597.4]
  assign regs_140_clock = clock; // @[:@135606.4]
  assign regs_140_reset = io_reset; // @[:@135607.4 RegFile.scala 76:16:@135614.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@135613.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@135617.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@135611.4]
  assign regs_141_clock = clock; // @[:@135620.4]
  assign regs_141_reset = io_reset; // @[:@135621.4 RegFile.scala 76:16:@135628.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@135627.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@135631.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@135625.4]
  assign regs_142_clock = clock; // @[:@135634.4]
  assign regs_142_reset = io_reset; // @[:@135635.4 RegFile.scala 76:16:@135642.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@135641.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@135645.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@135639.4]
  assign regs_143_clock = clock; // @[:@135648.4]
  assign regs_143_reset = io_reset; // @[:@135649.4 RegFile.scala 76:16:@135656.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@135655.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@135659.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@135653.4]
  assign regs_144_clock = clock; // @[:@135662.4]
  assign regs_144_reset = io_reset; // @[:@135663.4 RegFile.scala 76:16:@135670.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@135669.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@135673.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@135667.4]
  assign regs_145_clock = clock; // @[:@135676.4]
  assign regs_145_reset = io_reset; // @[:@135677.4 RegFile.scala 76:16:@135684.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@135683.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@135687.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@135681.4]
  assign regs_146_clock = clock; // @[:@135690.4]
  assign regs_146_reset = io_reset; // @[:@135691.4 RegFile.scala 76:16:@135698.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@135697.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@135701.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@135695.4]
  assign regs_147_clock = clock; // @[:@135704.4]
  assign regs_147_reset = io_reset; // @[:@135705.4 RegFile.scala 76:16:@135712.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@135711.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@135715.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@135709.4]
  assign regs_148_clock = clock; // @[:@135718.4]
  assign regs_148_reset = io_reset; // @[:@135719.4 RegFile.scala 76:16:@135726.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@135725.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@135729.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@135723.4]
  assign regs_149_clock = clock; // @[:@135732.4]
  assign regs_149_reset = io_reset; // @[:@135733.4 RegFile.scala 76:16:@135740.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@135739.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@135743.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@135737.4]
  assign regs_150_clock = clock; // @[:@135746.4]
  assign regs_150_reset = io_reset; // @[:@135747.4 RegFile.scala 76:16:@135754.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@135753.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@135757.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@135751.4]
  assign regs_151_clock = clock; // @[:@135760.4]
  assign regs_151_reset = io_reset; // @[:@135761.4 RegFile.scala 76:16:@135768.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@135767.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@135771.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@135765.4]
  assign regs_152_clock = clock; // @[:@135774.4]
  assign regs_152_reset = io_reset; // @[:@135775.4 RegFile.scala 76:16:@135782.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@135781.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@135785.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@135779.4]
  assign regs_153_clock = clock; // @[:@135788.4]
  assign regs_153_reset = io_reset; // @[:@135789.4 RegFile.scala 76:16:@135796.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@135795.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@135799.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@135793.4]
  assign regs_154_clock = clock; // @[:@135802.4]
  assign regs_154_reset = io_reset; // @[:@135803.4 RegFile.scala 76:16:@135810.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@135809.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@135813.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@135807.4]
  assign regs_155_clock = clock; // @[:@135816.4]
  assign regs_155_reset = io_reset; // @[:@135817.4 RegFile.scala 76:16:@135824.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@135823.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@135827.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@135821.4]
  assign regs_156_clock = clock; // @[:@135830.4]
  assign regs_156_reset = io_reset; // @[:@135831.4 RegFile.scala 76:16:@135838.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@135837.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@135841.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@135835.4]
  assign regs_157_clock = clock; // @[:@135844.4]
  assign regs_157_reset = io_reset; // @[:@135845.4 RegFile.scala 76:16:@135852.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@135851.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@135855.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@135849.4]
  assign regs_158_clock = clock; // @[:@135858.4]
  assign regs_158_reset = io_reset; // @[:@135859.4 RegFile.scala 76:16:@135866.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@135865.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@135869.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@135863.4]
  assign regs_159_clock = clock; // @[:@135872.4]
  assign regs_159_reset = io_reset; // @[:@135873.4 RegFile.scala 76:16:@135880.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@135879.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@135883.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@135877.4]
  assign regs_160_clock = clock; // @[:@135886.4]
  assign regs_160_reset = io_reset; // @[:@135887.4 RegFile.scala 76:16:@135894.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@135893.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@135897.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@135891.4]
  assign regs_161_clock = clock; // @[:@135900.4]
  assign regs_161_reset = io_reset; // @[:@135901.4 RegFile.scala 76:16:@135908.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@135907.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@135911.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@135905.4]
  assign regs_162_clock = clock; // @[:@135914.4]
  assign regs_162_reset = io_reset; // @[:@135915.4 RegFile.scala 76:16:@135922.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@135921.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@135925.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@135919.4]
  assign regs_163_clock = clock; // @[:@135928.4]
  assign regs_163_reset = io_reset; // @[:@135929.4 RegFile.scala 76:16:@135936.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@135935.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@135939.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@135933.4]
  assign regs_164_clock = clock; // @[:@135942.4]
  assign regs_164_reset = io_reset; // @[:@135943.4 RegFile.scala 76:16:@135950.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@135949.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@135953.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@135947.4]
  assign regs_165_clock = clock; // @[:@135956.4]
  assign regs_165_reset = io_reset; // @[:@135957.4 RegFile.scala 76:16:@135964.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@135963.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@135967.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@135961.4]
  assign regs_166_clock = clock; // @[:@135970.4]
  assign regs_166_reset = io_reset; // @[:@135971.4 RegFile.scala 76:16:@135978.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@135977.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@135981.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@135975.4]
  assign regs_167_clock = clock; // @[:@135984.4]
  assign regs_167_reset = io_reset; // @[:@135985.4 RegFile.scala 76:16:@135992.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@135991.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@135995.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@135989.4]
  assign regs_168_clock = clock; // @[:@135998.4]
  assign regs_168_reset = io_reset; // @[:@135999.4 RegFile.scala 76:16:@136006.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@136005.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@136009.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@136003.4]
  assign regs_169_clock = clock; // @[:@136012.4]
  assign regs_169_reset = io_reset; // @[:@136013.4 RegFile.scala 76:16:@136020.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@136019.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@136023.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@136017.4]
  assign regs_170_clock = clock; // @[:@136026.4]
  assign regs_170_reset = io_reset; // @[:@136027.4 RegFile.scala 76:16:@136034.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@136033.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@136037.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@136031.4]
  assign regs_171_clock = clock; // @[:@136040.4]
  assign regs_171_reset = io_reset; // @[:@136041.4 RegFile.scala 76:16:@136048.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@136047.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@136051.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@136045.4]
  assign regs_172_clock = clock; // @[:@136054.4]
  assign regs_172_reset = io_reset; // @[:@136055.4 RegFile.scala 76:16:@136062.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@136061.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@136065.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@136059.4]
  assign regs_173_clock = clock; // @[:@136068.4]
  assign regs_173_reset = io_reset; // @[:@136069.4 RegFile.scala 76:16:@136076.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@136075.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@136079.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@136073.4]
  assign regs_174_clock = clock; // @[:@136082.4]
  assign regs_174_reset = io_reset; // @[:@136083.4 RegFile.scala 76:16:@136090.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@136089.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@136093.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@136087.4]
  assign regs_175_clock = clock; // @[:@136096.4]
  assign regs_175_reset = io_reset; // @[:@136097.4 RegFile.scala 76:16:@136104.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@136103.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@136107.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@136101.4]
  assign regs_176_clock = clock; // @[:@136110.4]
  assign regs_176_reset = io_reset; // @[:@136111.4 RegFile.scala 76:16:@136118.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@136117.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@136121.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@136115.4]
  assign regs_177_clock = clock; // @[:@136124.4]
  assign regs_177_reset = io_reset; // @[:@136125.4 RegFile.scala 76:16:@136132.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@136131.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@136135.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@136129.4]
  assign regs_178_clock = clock; // @[:@136138.4]
  assign regs_178_reset = io_reset; // @[:@136139.4 RegFile.scala 76:16:@136146.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@136145.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@136149.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@136143.4]
  assign regs_179_clock = clock; // @[:@136152.4]
  assign regs_179_reset = io_reset; // @[:@136153.4 RegFile.scala 76:16:@136160.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@136159.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@136163.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@136157.4]
  assign regs_180_clock = clock; // @[:@136166.4]
  assign regs_180_reset = io_reset; // @[:@136167.4 RegFile.scala 76:16:@136174.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@136173.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@136177.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@136171.4]
  assign regs_181_clock = clock; // @[:@136180.4]
  assign regs_181_reset = io_reset; // @[:@136181.4 RegFile.scala 76:16:@136188.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@136187.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@136191.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@136185.4]
  assign regs_182_clock = clock; // @[:@136194.4]
  assign regs_182_reset = io_reset; // @[:@136195.4 RegFile.scala 76:16:@136202.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@136201.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@136205.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@136199.4]
  assign regs_183_clock = clock; // @[:@136208.4]
  assign regs_183_reset = io_reset; // @[:@136209.4 RegFile.scala 76:16:@136216.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@136215.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@136219.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@136213.4]
  assign regs_184_clock = clock; // @[:@136222.4]
  assign regs_184_reset = io_reset; // @[:@136223.4 RegFile.scala 76:16:@136230.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@136229.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@136233.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@136227.4]
  assign regs_185_clock = clock; // @[:@136236.4]
  assign regs_185_reset = io_reset; // @[:@136237.4 RegFile.scala 76:16:@136244.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@136243.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@136247.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@136241.4]
  assign regs_186_clock = clock; // @[:@136250.4]
  assign regs_186_reset = io_reset; // @[:@136251.4 RegFile.scala 76:16:@136258.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@136257.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@136261.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@136255.4]
  assign regs_187_clock = clock; // @[:@136264.4]
  assign regs_187_reset = io_reset; // @[:@136265.4 RegFile.scala 76:16:@136272.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@136271.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@136275.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@136269.4]
  assign regs_188_clock = clock; // @[:@136278.4]
  assign regs_188_reset = io_reset; // @[:@136279.4 RegFile.scala 76:16:@136286.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@136285.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@136289.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@136283.4]
  assign regs_189_clock = clock; // @[:@136292.4]
  assign regs_189_reset = io_reset; // @[:@136293.4 RegFile.scala 76:16:@136300.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@136299.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@136303.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@136297.4]
  assign regs_190_clock = clock; // @[:@136306.4]
  assign regs_190_reset = io_reset; // @[:@136307.4 RegFile.scala 76:16:@136314.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@136313.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@136317.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@136311.4]
  assign regs_191_clock = clock; // @[:@136320.4]
  assign regs_191_reset = io_reset; // @[:@136321.4 RegFile.scala 76:16:@136328.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@136327.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@136331.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@136325.4]
  assign regs_192_clock = clock; // @[:@136334.4]
  assign regs_192_reset = io_reset; // @[:@136335.4 RegFile.scala 76:16:@136342.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@136341.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@136345.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@136339.4]
  assign regs_193_clock = clock; // @[:@136348.4]
  assign regs_193_reset = io_reset; // @[:@136349.4 RegFile.scala 76:16:@136356.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@136355.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@136359.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@136353.4]
  assign regs_194_clock = clock; // @[:@136362.4]
  assign regs_194_reset = io_reset; // @[:@136363.4 RegFile.scala 76:16:@136370.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@136369.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@136373.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@136367.4]
  assign regs_195_clock = clock; // @[:@136376.4]
  assign regs_195_reset = io_reset; // @[:@136377.4 RegFile.scala 76:16:@136384.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@136383.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@136387.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@136381.4]
  assign regs_196_clock = clock; // @[:@136390.4]
  assign regs_196_reset = io_reset; // @[:@136391.4 RegFile.scala 76:16:@136398.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@136397.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@136401.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@136395.4]
  assign regs_197_clock = clock; // @[:@136404.4]
  assign regs_197_reset = io_reset; // @[:@136405.4 RegFile.scala 76:16:@136412.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@136411.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@136415.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@136409.4]
  assign regs_198_clock = clock; // @[:@136418.4]
  assign regs_198_reset = io_reset; // @[:@136419.4 RegFile.scala 76:16:@136426.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@136425.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@136429.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@136423.4]
  assign regs_199_clock = clock; // @[:@136432.4]
  assign regs_199_reset = io_reset; // @[:@136433.4 RegFile.scala 76:16:@136440.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@136439.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@136443.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@136437.4]
  assign regs_200_clock = clock; // @[:@136446.4]
  assign regs_200_reset = io_reset; // @[:@136447.4 RegFile.scala 76:16:@136454.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@136453.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@136457.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@136451.4]
  assign regs_201_clock = clock; // @[:@136460.4]
  assign regs_201_reset = io_reset; // @[:@136461.4 RegFile.scala 76:16:@136468.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@136467.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@136471.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@136465.4]
  assign regs_202_clock = clock; // @[:@136474.4]
  assign regs_202_reset = io_reset; // @[:@136475.4 RegFile.scala 76:16:@136482.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@136481.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@136485.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@136479.4]
  assign regs_203_clock = clock; // @[:@136488.4]
  assign regs_203_reset = io_reset; // @[:@136489.4 RegFile.scala 76:16:@136496.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@136495.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@136499.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@136493.4]
  assign regs_204_clock = clock; // @[:@136502.4]
  assign regs_204_reset = io_reset; // @[:@136503.4 RegFile.scala 76:16:@136510.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@136509.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@136513.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@136507.4]
  assign regs_205_clock = clock; // @[:@136516.4]
  assign regs_205_reset = io_reset; // @[:@136517.4 RegFile.scala 76:16:@136524.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@136523.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@136527.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@136521.4]
  assign regs_206_clock = clock; // @[:@136530.4]
  assign regs_206_reset = io_reset; // @[:@136531.4 RegFile.scala 76:16:@136538.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@136537.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@136541.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@136535.4]
  assign regs_207_clock = clock; // @[:@136544.4]
  assign regs_207_reset = io_reset; // @[:@136545.4 RegFile.scala 76:16:@136552.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@136551.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@136555.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@136549.4]
  assign regs_208_clock = clock; // @[:@136558.4]
  assign regs_208_reset = io_reset; // @[:@136559.4 RegFile.scala 76:16:@136566.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@136565.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@136569.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@136563.4]
  assign regs_209_clock = clock; // @[:@136572.4]
  assign regs_209_reset = io_reset; // @[:@136573.4 RegFile.scala 76:16:@136580.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@136579.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@136583.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@136577.4]
  assign regs_210_clock = clock; // @[:@136586.4]
  assign regs_210_reset = io_reset; // @[:@136587.4 RegFile.scala 76:16:@136594.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@136593.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@136597.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@136591.4]
  assign regs_211_clock = clock; // @[:@136600.4]
  assign regs_211_reset = io_reset; // @[:@136601.4 RegFile.scala 76:16:@136608.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@136607.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@136611.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@136605.4]
  assign regs_212_clock = clock; // @[:@136614.4]
  assign regs_212_reset = io_reset; // @[:@136615.4 RegFile.scala 76:16:@136622.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@136621.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@136625.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@136619.4]
  assign regs_213_clock = clock; // @[:@136628.4]
  assign regs_213_reset = io_reset; // @[:@136629.4 RegFile.scala 76:16:@136636.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@136635.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@136639.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@136633.4]
  assign regs_214_clock = clock; // @[:@136642.4]
  assign regs_214_reset = io_reset; // @[:@136643.4 RegFile.scala 76:16:@136650.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@136649.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@136653.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@136647.4]
  assign regs_215_clock = clock; // @[:@136656.4]
  assign regs_215_reset = io_reset; // @[:@136657.4 RegFile.scala 76:16:@136664.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@136663.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@136667.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@136661.4]
  assign regs_216_clock = clock; // @[:@136670.4]
  assign regs_216_reset = io_reset; // @[:@136671.4 RegFile.scala 76:16:@136678.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@136677.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@136681.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@136675.4]
  assign regs_217_clock = clock; // @[:@136684.4]
  assign regs_217_reset = io_reset; // @[:@136685.4 RegFile.scala 76:16:@136692.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@136691.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@136695.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@136689.4]
  assign regs_218_clock = clock; // @[:@136698.4]
  assign regs_218_reset = io_reset; // @[:@136699.4 RegFile.scala 76:16:@136706.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@136705.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@136709.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@136703.4]
  assign regs_219_clock = clock; // @[:@136712.4]
  assign regs_219_reset = io_reset; // @[:@136713.4 RegFile.scala 76:16:@136720.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@136719.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@136723.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@136717.4]
  assign regs_220_clock = clock; // @[:@136726.4]
  assign regs_220_reset = io_reset; // @[:@136727.4 RegFile.scala 76:16:@136734.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@136733.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@136737.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@136731.4]
  assign regs_221_clock = clock; // @[:@136740.4]
  assign regs_221_reset = io_reset; // @[:@136741.4 RegFile.scala 76:16:@136748.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@136747.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@136751.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@136745.4]
  assign regs_222_clock = clock; // @[:@136754.4]
  assign regs_222_reset = io_reset; // @[:@136755.4 RegFile.scala 76:16:@136762.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@136761.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@136765.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@136759.4]
  assign regs_223_clock = clock; // @[:@136768.4]
  assign regs_223_reset = io_reset; // @[:@136769.4 RegFile.scala 76:16:@136776.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@136775.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@136779.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@136773.4]
  assign regs_224_clock = clock; // @[:@136782.4]
  assign regs_224_reset = io_reset; // @[:@136783.4 RegFile.scala 76:16:@136790.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@136789.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@136793.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@136787.4]
  assign regs_225_clock = clock; // @[:@136796.4]
  assign regs_225_reset = io_reset; // @[:@136797.4 RegFile.scala 76:16:@136804.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@136803.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@136807.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@136801.4]
  assign regs_226_clock = clock; // @[:@136810.4]
  assign regs_226_reset = io_reset; // @[:@136811.4 RegFile.scala 76:16:@136818.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@136817.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@136821.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@136815.4]
  assign regs_227_clock = clock; // @[:@136824.4]
  assign regs_227_reset = io_reset; // @[:@136825.4 RegFile.scala 76:16:@136832.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@136831.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@136835.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@136829.4]
  assign regs_228_clock = clock; // @[:@136838.4]
  assign regs_228_reset = io_reset; // @[:@136839.4 RegFile.scala 76:16:@136846.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@136845.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@136849.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@136843.4]
  assign regs_229_clock = clock; // @[:@136852.4]
  assign regs_229_reset = io_reset; // @[:@136853.4 RegFile.scala 76:16:@136860.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@136859.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@136863.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@136857.4]
  assign regs_230_clock = clock; // @[:@136866.4]
  assign regs_230_reset = io_reset; // @[:@136867.4 RegFile.scala 76:16:@136874.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@136873.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@136877.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@136871.4]
  assign regs_231_clock = clock; // @[:@136880.4]
  assign regs_231_reset = io_reset; // @[:@136881.4 RegFile.scala 76:16:@136888.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@136887.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@136891.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@136885.4]
  assign regs_232_clock = clock; // @[:@136894.4]
  assign regs_232_reset = io_reset; // @[:@136895.4 RegFile.scala 76:16:@136902.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@136901.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@136905.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@136899.4]
  assign regs_233_clock = clock; // @[:@136908.4]
  assign regs_233_reset = io_reset; // @[:@136909.4 RegFile.scala 76:16:@136916.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@136915.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@136919.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@136913.4]
  assign regs_234_clock = clock; // @[:@136922.4]
  assign regs_234_reset = io_reset; // @[:@136923.4 RegFile.scala 76:16:@136930.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@136929.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@136933.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@136927.4]
  assign regs_235_clock = clock; // @[:@136936.4]
  assign regs_235_reset = io_reset; // @[:@136937.4 RegFile.scala 76:16:@136944.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@136943.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@136947.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@136941.4]
  assign regs_236_clock = clock; // @[:@136950.4]
  assign regs_236_reset = io_reset; // @[:@136951.4 RegFile.scala 76:16:@136958.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@136957.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@136961.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@136955.4]
  assign regs_237_clock = clock; // @[:@136964.4]
  assign regs_237_reset = io_reset; // @[:@136965.4 RegFile.scala 76:16:@136972.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@136971.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@136975.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@136969.4]
  assign regs_238_clock = clock; // @[:@136978.4]
  assign regs_238_reset = io_reset; // @[:@136979.4 RegFile.scala 76:16:@136986.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@136985.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@136989.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@136983.4]
  assign regs_239_clock = clock; // @[:@136992.4]
  assign regs_239_reset = io_reset; // @[:@136993.4 RegFile.scala 76:16:@137000.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@136999.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@137003.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@136997.4]
  assign regs_240_clock = clock; // @[:@137006.4]
  assign regs_240_reset = io_reset; // @[:@137007.4 RegFile.scala 76:16:@137014.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@137013.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@137017.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@137011.4]
  assign regs_241_clock = clock; // @[:@137020.4]
  assign regs_241_reset = io_reset; // @[:@137021.4 RegFile.scala 76:16:@137028.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@137027.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@137031.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@137025.4]
  assign regs_242_clock = clock; // @[:@137034.4]
  assign regs_242_reset = io_reset; // @[:@137035.4 RegFile.scala 76:16:@137042.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@137041.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@137045.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@137039.4]
  assign regs_243_clock = clock; // @[:@137048.4]
  assign regs_243_reset = io_reset; // @[:@137049.4 RegFile.scala 76:16:@137056.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@137055.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@137059.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@137053.4]
  assign regs_244_clock = clock; // @[:@137062.4]
  assign regs_244_reset = io_reset; // @[:@137063.4 RegFile.scala 76:16:@137070.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@137069.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@137073.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@137067.4]
  assign regs_245_clock = clock; // @[:@137076.4]
  assign regs_245_reset = io_reset; // @[:@137077.4 RegFile.scala 76:16:@137084.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@137083.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@137087.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@137081.4]
  assign regs_246_clock = clock; // @[:@137090.4]
  assign regs_246_reset = io_reset; // @[:@137091.4 RegFile.scala 76:16:@137098.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@137097.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@137101.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@137095.4]
  assign regs_247_clock = clock; // @[:@137104.4]
  assign regs_247_reset = io_reset; // @[:@137105.4 RegFile.scala 76:16:@137112.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@137111.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@137115.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@137109.4]
  assign regs_248_clock = clock; // @[:@137118.4]
  assign regs_248_reset = io_reset; // @[:@137119.4 RegFile.scala 76:16:@137126.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@137125.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@137129.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@137123.4]
  assign regs_249_clock = clock; // @[:@137132.4]
  assign regs_249_reset = io_reset; // @[:@137133.4 RegFile.scala 76:16:@137140.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@137139.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@137143.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@137137.4]
  assign regs_250_clock = clock; // @[:@137146.4]
  assign regs_250_reset = io_reset; // @[:@137147.4 RegFile.scala 76:16:@137154.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@137153.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@137157.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@137151.4]
  assign regs_251_clock = clock; // @[:@137160.4]
  assign regs_251_reset = io_reset; // @[:@137161.4 RegFile.scala 76:16:@137168.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@137167.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@137171.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@137165.4]
  assign regs_252_clock = clock; // @[:@137174.4]
  assign regs_252_reset = io_reset; // @[:@137175.4 RegFile.scala 76:16:@137182.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@137181.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@137185.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@137179.4]
  assign regs_253_clock = clock; // @[:@137188.4]
  assign regs_253_reset = io_reset; // @[:@137189.4 RegFile.scala 76:16:@137196.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@137195.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@137199.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@137193.4]
  assign regs_254_clock = clock; // @[:@137202.4]
  assign regs_254_reset = io_reset; // @[:@137203.4 RegFile.scala 76:16:@137210.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@137209.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@137213.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@137207.4]
  assign regs_255_clock = clock; // @[:@137216.4]
  assign regs_255_reset = io_reset; // @[:@137217.4 RegFile.scala 76:16:@137224.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@137223.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@137227.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@137221.4]
  assign regs_256_clock = clock; // @[:@137230.4]
  assign regs_256_reset = io_reset; // @[:@137231.4 RegFile.scala 76:16:@137238.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@137237.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@137241.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@137235.4]
  assign regs_257_clock = clock; // @[:@137244.4]
  assign regs_257_reset = io_reset; // @[:@137245.4 RegFile.scala 76:16:@137252.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@137251.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@137255.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@137249.4]
  assign regs_258_clock = clock; // @[:@137258.4]
  assign regs_258_reset = io_reset; // @[:@137259.4 RegFile.scala 76:16:@137266.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@137265.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@137269.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@137263.4]
  assign regs_259_clock = clock; // @[:@137272.4]
  assign regs_259_reset = io_reset; // @[:@137273.4 RegFile.scala 76:16:@137280.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@137279.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@137283.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@137277.4]
  assign regs_260_clock = clock; // @[:@137286.4]
  assign regs_260_reset = io_reset; // @[:@137287.4 RegFile.scala 76:16:@137294.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@137293.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@137297.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@137291.4]
  assign regs_261_clock = clock; // @[:@137300.4]
  assign regs_261_reset = io_reset; // @[:@137301.4 RegFile.scala 76:16:@137308.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@137307.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@137311.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@137305.4]
  assign regs_262_clock = clock; // @[:@137314.4]
  assign regs_262_reset = io_reset; // @[:@137315.4 RegFile.scala 76:16:@137322.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@137321.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@137325.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@137319.4]
  assign regs_263_clock = clock; // @[:@137328.4]
  assign regs_263_reset = io_reset; // @[:@137329.4 RegFile.scala 76:16:@137336.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@137335.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@137339.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@137333.4]
  assign regs_264_clock = clock; // @[:@137342.4]
  assign regs_264_reset = io_reset; // @[:@137343.4 RegFile.scala 76:16:@137350.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@137349.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@137353.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@137347.4]
  assign regs_265_clock = clock; // @[:@137356.4]
  assign regs_265_reset = io_reset; // @[:@137357.4 RegFile.scala 76:16:@137364.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@137363.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@137367.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@137361.4]
  assign regs_266_clock = clock; // @[:@137370.4]
  assign regs_266_reset = io_reset; // @[:@137371.4 RegFile.scala 76:16:@137378.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@137377.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@137381.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@137375.4]
  assign regs_267_clock = clock; // @[:@137384.4]
  assign regs_267_reset = io_reset; // @[:@137385.4 RegFile.scala 76:16:@137392.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@137391.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@137395.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@137389.4]
  assign regs_268_clock = clock; // @[:@137398.4]
  assign regs_268_reset = io_reset; // @[:@137399.4 RegFile.scala 76:16:@137406.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@137405.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@137409.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@137403.4]
  assign regs_269_clock = clock; // @[:@137412.4]
  assign regs_269_reset = io_reset; // @[:@137413.4 RegFile.scala 76:16:@137420.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@137419.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@137423.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@137417.4]
  assign regs_270_clock = clock; // @[:@137426.4]
  assign regs_270_reset = io_reset; // @[:@137427.4 RegFile.scala 76:16:@137434.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@137433.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@137437.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@137431.4]
  assign regs_271_clock = clock; // @[:@137440.4]
  assign regs_271_reset = io_reset; // @[:@137441.4 RegFile.scala 76:16:@137448.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@137447.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@137451.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@137445.4]
  assign regs_272_clock = clock; // @[:@137454.4]
  assign regs_272_reset = io_reset; // @[:@137455.4 RegFile.scala 76:16:@137462.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@137461.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@137465.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@137459.4]
  assign regs_273_clock = clock; // @[:@137468.4]
  assign regs_273_reset = io_reset; // @[:@137469.4 RegFile.scala 76:16:@137476.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@137475.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@137479.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@137473.4]
  assign regs_274_clock = clock; // @[:@137482.4]
  assign regs_274_reset = io_reset; // @[:@137483.4 RegFile.scala 76:16:@137490.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@137489.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@137493.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@137487.4]
  assign regs_275_clock = clock; // @[:@137496.4]
  assign regs_275_reset = io_reset; // @[:@137497.4 RegFile.scala 76:16:@137504.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@137503.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@137507.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@137501.4]
  assign regs_276_clock = clock; // @[:@137510.4]
  assign regs_276_reset = io_reset; // @[:@137511.4 RegFile.scala 76:16:@137518.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@137517.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@137521.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@137515.4]
  assign regs_277_clock = clock; // @[:@137524.4]
  assign regs_277_reset = io_reset; // @[:@137525.4 RegFile.scala 76:16:@137532.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@137531.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@137535.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@137529.4]
  assign regs_278_clock = clock; // @[:@137538.4]
  assign regs_278_reset = io_reset; // @[:@137539.4 RegFile.scala 76:16:@137546.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@137545.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@137549.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@137543.4]
  assign regs_279_clock = clock; // @[:@137552.4]
  assign regs_279_reset = io_reset; // @[:@137553.4 RegFile.scala 76:16:@137560.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@137559.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@137563.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@137557.4]
  assign regs_280_clock = clock; // @[:@137566.4]
  assign regs_280_reset = io_reset; // @[:@137567.4 RegFile.scala 76:16:@137574.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@137573.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@137577.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@137571.4]
  assign regs_281_clock = clock; // @[:@137580.4]
  assign regs_281_reset = io_reset; // @[:@137581.4 RegFile.scala 76:16:@137588.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@137587.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@137591.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@137585.4]
  assign regs_282_clock = clock; // @[:@137594.4]
  assign regs_282_reset = io_reset; // @[:@137595.4 RegFile.scala 76:16:@137602.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@137601.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@137605.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@137599.4]
  assign regs_283_clock = clock; // @[:@137608.4]
  assign regs_283_reset = io_reset; // @[:@137609.4 RegFile.scala 76:16:@137616.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@137615.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@137619.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@137613.4]
  assign regs_284_clock = clock; // @[:@137622.4]
  assign regs_284_reset = io_reset; // @[:@137623.4 RegFile.scala 76:16:@137630.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@137629.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@137633.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@137627.4]
  assign regs_285_clock = clock; // @[:@137636.4]
  assign regs_285_reset = io_reset; // @[:@137637.4 RegFile.scala 76:16:@137644.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@137643.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@137647.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@137641.4]
  assign regs_286_clock = clock; // @[:@137650.4]
  assign regs_286_reset = io_reset; // @[:@137651.4 RegFile.scala 76:16:@137658.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@137657.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@137661.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@137655.4]
  assign regs_287_clock = clock; // @[:@137664.4]
  assign regs_287_reset = io_reset; // @[:@137665.4 RegFile.scala 76:16:@137672.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@137671.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@137675.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@137669.4]
  assign regs_288_clock = clock; // @[:@137678.4]
  assign regs_288_reset = io_reset; // @[:@137679.4 RegFile.scala 76:16:@137686.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@137685.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@137689.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@137683.4]
  assign regs_289_clock = clock; // @[:@137692.4]
  assign regs_289_reset = io_reset; // @[:@137693.4 RegFile.scala 76:16:@137700.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@137699.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@137703.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@137697.4]
  assign regs_290_clock = clock; // @[:@137706.4]
  assign regs_290_reset = io_reset; // @[:@137707.4 RegFile.scala 76:16:@137714.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@137713.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@137717.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@137711.4]
  assign regs_291_clock = clock; // @[:@137720.4]
  assign regs_291_reset = io_reset; // @[:@137721.4 RegFile.scala 76:16:@137728.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@137727.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@137731.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@137725.4]
  assign regs_292_clock = clock; // @[:@137734.4]
  assign regs_292_reset = io_reset; // @[:@137735.4 RegFile.scala 76:16:@137742.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@137741.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@137745.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@137739.4]
  assign regs_293_clock = clock; // @[:@137748.4]
  assign regs_293_reset = io_reset; // @[:@137749.4 RegFile.scala 76:16:@137756.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@137755.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@137759.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@137753.4]
  assign regs_294_clock = clock; // @[:@137762.4]
  assign regs_294_reset = io_reset; // @[:@137763.4 RegFile.scala 76:16:@137770.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@137769.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@137773.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@137767.4]
  assign regs_295_clock = clock; // @[:@137776.4]
  assign regs_295_reset = io_reset; // @[:@137777.4 RegFile.scala 76:16:@137784.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@137783.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@137787.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@137781.4]
  assign regs_296_clock = clock; // @[:@137790.4]
  assign regs_296_reset = io_reset; // @[:@137791.4 RegFile.scala 76:16:@137798.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@137797.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@137801.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@137795.4]
  assign regs_297_clock = clock; // @[:@137804.4]
  assign regs_297_reset = io_reset; // @[:@137805.4 RegFile.scala 76:16:@137812.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@137811.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@137815.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@137809.4]
  assign regs_298_clock = clock; // @[:@137818.4]
  assign regs_298_reset = io_reset; // @[:@137819.4 RegFile.scala 76:16:@137826.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@137825.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@137829.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@137823.4]
  assign regs_299_clock = clock; // @[:@137832.4]
  assign regs_299_reset = io_reset; // @[:@137833.4 RegFile.scala 76:16:@137840.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@137839.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@137843.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@137837.4]
  assign regs_300_clock = clock; // @[:@137846.4]
  assign regs_300_reset = io_reset; // @[:@137847.4 RegFile.scala 76:16:@137854.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@137853.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@137857.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@137851.4]
  assign regs_301_clock = clock; // @[:@137860.4]
  assign regs_301_reset = io_reset; // @[:@137861.4 RegFile.scala 76:16:@137868.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@137867.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@137871.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@137865.4]
  assign regs_302_clock = clock; // @[:@137874.4]
  assign regs_302_reset = io_reset; // @[:@137875.4 RegFile.scala 76:16:@137882.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@137881.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@137885.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@137879.4]
  assign regs_303_clock = clock; // @[:@137888.4]
  assign regs_303_reset = io_reset; // @[:@137889.4 RegFile.scala 76:16:@137896.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@137895.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@137899.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@137893.4]
  assign regs_304_clock = clock; // @[:@137902.4]
  assign regs_304_reset = io_reset; // @[:@137903.4 RegFile.scala 76:16:@137910.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@137909.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@137913.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@137907.4]
  assign regs_305_clock = clock; // @[:@137916.4]
  assign regs_305_reset = io_reset; // @[:@137917.4 RegFile.scala 76:16:@137924.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@137923.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@137927.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@137921.4]
  assign regs_306_clock = clock; // @[:@137930.4]
  assign regs_306_reset = io_reset; // @[:@137931.4 RegFile.scala 76:16:@137938.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@137937.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@137941.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@137935.4]
  assign regs_307_clock = clock; // @[:@137944.4]
  assign regs_307_reset = io_reset; // @[:@137945.4 RegFile.scala 76:16:@137952.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@137951.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@137955.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@137949.4]
  assign regs_308_clock = clock; // @[:@137958.4]
  assign regs_308_reset = io_reset; // @[:@137959.4 RegFile.scala 76:16:@137966.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@137965.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@137969.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@137963.4]
  assign regs_309_clock = clock; // @[:@137972.4]
  assign regs_309_reset = io_reset; // @[:@137973.4 RegFile.scala 76:16:@137980.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@137979.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@137983.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@137977.4]
  assign regs_310_clock = clock; // @[:@137986.4]
  assign regs_310_reset = io_reset; // @[:@137987.4 RegFile.scala 76:16:@137994.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@137993.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@137997.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@137991.4]
  assign regs_311_clock = clock; // @[:@138000.4]
  assign regs_311_reset = io_reset; // @[:@138001.4 RegFile.scala 76:16:@138008.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@138007.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@138011.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@138005.4]
  assign regs_312_clock = clock; // @[:@138014.4]
  assign regs_312_reset = io_reset; // @[:@138015.4 RegFile.scala 76:16:@138022.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@138021.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@138025.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@138019.4]
  assign regs_313_clock = clock; // @[:@138028.4]
  assign regs_313_reset = io_reset; // @[:@138029.4 RegFile.scala 76:16:@138036.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@138035.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@138039.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@138033.4]
  assign regs_314_clock = clock; // @[:@138042.4]
  assign regs_314_reset = io_reset; // @[:@138043.4 RegFile.scala 76:16:@138050.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@138049.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@138053.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@138047.4]
  assign regs_315_clock = clock; // @[:@138056.4]
  assign regs_315_reset = io_reset; // @[:@138057.4 RegFile.scala 76:16:@138064.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@138063.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@138067.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@138061.4]
  assign regs_316_clock = clock; // @[:@138070.4]
  assign regs_316_reset = io_reset; // @[:@138071.4 RegFile.scala 76:16:@138078.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@138077.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@138081.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@138075.4]
  assign regs_317_clock = clock; // @[:@138084.4]
  assign regs_317_reset = io_reset; // @[:@138085.4 RegFile.scala 76:16:@138092.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@138091.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@138095.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@138089.4]
  assign regs_318_clock = clock; // @[:@138098.4]
  assign regs_318_reset = io_reset; // @[:@138099.4 RegFile.scala 76:16:@138106.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@138105.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@138109.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@138103.4]
  assign regs_319_clock = clock; // @[:@138112.4]
  assign regs_319_reset = io_reset; // @[:@138113.4 RegFile.scala 76:16:@138120.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@138119.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@138123.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@138117.4]
  assign regs_320_clock = clock; // @[:@138126.4]
  assign regs_320_reset = io_reset; // @[:@138127.4 RegFile.scala 76:16:@138134.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@138133.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@138137.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@138131.4]
  assign regs_321_clock = clock; // @[:@138140.4]
  assign regs_321_reset = io_reset; // @[:@138141.4 RegFile.scala 76:16:@138148.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@138147.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@138151.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@138145.4]
  assign regs_322_clock = clock; // @[:@138154.4]
  assign regs_322_reset = io_reset; // @[:@138155.4 RegFile.scala 76:16:@138162.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@138161.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@138165.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@138159.4]
  assign regs_323_clock = clock; // @[:@138168.4]
  assign regs_323_reset = io_reset; // @[:@138169.4 RegFile.scala 76:16:@138176.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@138175.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@138179.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@138173.4]
  assign regs_324_clock = clock; // @[:@138182.4]
  assign regs_324_reset = io_reset; // @[:@138183.4 RegFile.scala 76:16:@138190.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@138189.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@138193.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@138187.4]
  assign regs_325_clock = clock; // @[:@138196.4]
  assign regs_325_reset = io_reset; // @[:@138197.4 RegFile.scala 76:16:@138204.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@138203.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@138207.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@138201.4]
  assign regs_326_clock = clock; // @[:@138210.4]
  assign regs_326_reset = io_reset; // @[:@138211.4 RegFile.scala 76:16:@138218.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@138217.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@138221.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@138215.4]
  assign regs_327_clock = clock; // @[:@138224.4]
  assign regs_327_reset = io_reset; // @[:@138225.4 RegFile.scala 76:16:@138232.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@138231.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@138235.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@138229.4]
  assign regs_328_clock = clock; // @[:@138238.4]
  assign regs_328_reset = io_reset; // @[:@138239.4 RegFile.scala 76:16:@138246.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@138245.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@138249.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@138243.4]
  assign regs_329_clock = clock; // @[:@138252.4]
  assign regs_329_reset = io_reset; // @[:@138253.4 RegFile.scala 76:16:@138260.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@138259.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@138263.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@138257.4]
  assign regs_330_clock = clock; // @[:@138266.4]
  assign regs_330_reset = io_reset; // @[:@138267.4 RegFile.scala 76:16:@138274.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@138273.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@138277.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@138271.4]
  assign regs_331_clock = clock; // @[:@138280.4]
  assign regs_331_reset = io_reset; // @[:@138281.4 RegFile.scala 76:16:@138288.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@138287.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@138291.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@138285.4]
  assign regs_332_clock = clock; // @[:@138294.4]
  assign regs_332_reset = io_reset; // @[:@138295.4 RegFile.scala 76:16:@138302.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@138301.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@138305.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@138299.4]
  assign regs_333_clock = clock; // @[:@138308.4]
  assign regs_333_reset = io_reset; // @[:@138309.4 RegFile.scala 76:16:@138316.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@138315.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@138319.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@138313.4]
  assign regs_334_clock = clock; // @[:@138322.4]
  assign regs_334_reset = io_reset; // @[:@138323.4 RegFile.scala 76:16:@138330.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@138329.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@138333.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@138327.4]
  assign regs_335_clock = clock; // @[:@138336.4]
  assign regs_335_reset = io_reset; // @[:@138337.4 RegFile.scala 76:16:@138344.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@138343.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@138347.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@138341.4]
  assign regs_336_clock = clock; // @[:@138350.4]
  assign regs_336_reset = io_reset; // @[:@138351.4 RegFile.scala 76:16:@138358.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@138357.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@138361.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@138355.4]
  assign regs_337_clock = clock; // @[:@138364.4]
  assign regs_337_reset = io_reset; // @[:@138365.4 RegFile.scala 76:16:@138372.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@138371.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@138375.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@138369.4]
  assign regs_338_clock = clock; // @[:@138378.4]
  assign regs_338_reset = io_reset; // @[:@138379.4 RegFile.scala 76:16:@138386.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@138385.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@138389.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@138383.4]
  assign regs_339_clock = clock; // @[:@138392.4]
  assign regs_339_reset = io_reset; // @[:@138393.4 RegFile.scala 76:16:@138400.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@138399.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@138403.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@138397.4]
  assign regs_340_clock = clock; // @[:@138406.4]
  assign regs_340_reset = io_reset; // @[:@138407.4 RegFile.scala 76:16:@138414.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@138413.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@138417.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@138411.4]
  assign regs_341_clock = clock; // @[:@138420.4]
  assign regs_341_reset = io_reset; // @[:@138421.4 RegFile.scala 76:16:@138428.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@138427.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@138431.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@138425.4]
  assign regs_342_clock = clock; // @[:@138434.4]
  assign regs_342_reset = io_reset; // @[:@138435.4 RegFile.scala 76:16:@138442.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@138441.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@138445.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@138439.4]
  assign regs_343_clock = clock; // @[:@138448.4]
  assign regs_343_reset = io_reset; // @[:@138449.4 RegFile.scala 76:16:@138456.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@138455.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@138459.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@138453.4]
  assign regs_344_clock = clock; // @[:@138462.4]
  assign regs_344_reset = io_reset; // @[:@138463.4 RegFile.scala 76:16:@138470.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@138469.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@138473.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@138467.4]
  assign regs_345_clock = clock; // @[:@138476.4]
  assign regs_345_reset = io_reset; // @[:@138477.4 RegFile.scala 76:16:@138484.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@138483.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@138487.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@138481.4]
  assign regs_346_clock = clock; // @[:@138490.4]
  assign regs_346_reset = io_reset; // @[:@138491.4 RegFile.scala 76:16:@138498.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@138497.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@138501.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@138495.4]
  assign regs_347_clock = clock; // @[:@138504.4]
  assign regs_347_reset = io_reset; // @[:@138505.4 RegFile.scala 76:16:@138512.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@138511.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@138515.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@138509.4]
  assign regs_348_clock = clock; // @[:@138518.4]
  assign regs_348_reset = io_reset; // @[:@138519.4 RegFile.scala 76:16:@138526.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@138525.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@138529.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@138523.4]
  assign regs_349_clock = clock; // @[:@138532.4]
  assign regs_349_reset = io_reset; // @[:@138533.4 RegFile.scala 76:16:@138540.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@138539.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@138543.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@138537.4]
  assign regs_350_clock = clock; // @[:@138546.4]
  assign regs_350_reset = io_reset; // @[:@138547.4 RegFile.scala 76:16:@138554.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@138553.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@138557.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@138551.4]
  assign regs_351_clock = clock; // @[:@138560.4]
  assign regs_351_reset = io_reset; // @[:@138561.4 RegFile.scala 76:16:@138568.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@138567.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@138571.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@138565.4]
  assign regs_352_clock = clock; // @[:@138574.4]
  assign regs_352_reset = io_reset; // @[:@138575.4 RegFile.scala 76:16:@138582.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@138581.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@138585.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@138579.4]
  assign regs_353_clock = clock; // @[:@138588.4]
  assign regs_353_reset = io_reset; // @[:@138589.4 RegFile.scala 76:16:@138596.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@138595.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@138599.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@138593.4]
  assign regs_354_clock = clock; // @[:@138602.4]
  assign regs_354_reset = io_reset; // @[:@138603.4 RegFile.scala 76:16:@138610.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@138609.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@138613.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@138607.4]
  assign regs_355_clock = clock; // @[:@138616.4]
  assign regs_355_reset = io_reset; // @[:@138617.4 RegFile.scala 76:16:@138624.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@138623.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@138627.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@138621.4]
  assign regs_356_clock = clock; // @[:@138630.4]
  assign regs_356_reset = io_reset; // @[:@138631.4 RegFile.scala 76:16:@138638.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@138637.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@138641.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@138635.4]
  assign regs_357_clock = clock; // @[:@138644.4]
  assign regs_357_reset = io_reset; // @[:@138645.4 RegFile.scala 76:16:@138652.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@138651.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@138655.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@138649.4]
  assign regs_358_clock = clock; // @[:@138658.4]
  assign regs_358_reset = io_reset; // @[:@138659.4 RegFile.scala 76:16:@138666.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@138665.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@138669.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@138663.4]
  assign regs_359_clock = clock; // @[:@138672.4]
  assign regs_359_reset = io_reset; // @[:@138673.4 RegFile.scala 76:16:@138680.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@138679.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@138683.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@138677.4]
  assign regs_360_clock = clock; // @[:@138686.4]
  assign regs_360_reset = io_reset; // @[:@138687.4 RegFile.scala 76:16:@138694.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@138693.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@138697.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@138691.4]
  assign regs_361_clock = clock; // @[:@138700.4]
  assign regs_361_reset = io_reset; // @[:@138701.4 RegFile.scala 76:16:@138708.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@138707.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@138711.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@138705.4]
  assign regs_362_clock = clock; // @[:@138714.4]
  assign regs_362_reset = io_reset; // @[:@138715.4 RegFile.scala 76:16:@138722.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@138721.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@138725.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@138719.4]
  assign regs_363_clock = clock; // @[:@138728.4]
  assign regs_363_reset = io_reset; // @[:@138729.4 RegFile.scala 76:16:@138736.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@138735.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@138739.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@138733.4]
  assign regs_364_clock = clock; // @[:@138742.4]
  assign regs_364_reset = io_reset; // @[:@138743.4 RegFile.scala 76:16:@138750.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@138749.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@138753.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@138747.4]
  assign regs_365_clock = clock; // @[:@138756.4]
  assign regs_365_reset = io_reset; // @[:@138757.4 RegFile.scala 76:16:@138764.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@138763.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@138767.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@138761.4]
  assign regs_366_clock = clock; // @[:@138770.4]
  assign regs_366_reset = io_reset; // @[:@138771.4 RegFile.scala 76:16:@138778.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@138777.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@138781.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@138775.4]
  assign regs_367_clock = clock; // @[:@138784.4]
  assign regs_367_reset = io_reset; // @[:@138785.4 RegFile.scala 76:16:@138792.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@138791.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@138795.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@138789.4]
  assign regs_368_clock = clock; // @[:@138798.4]
  assign regs_368_reset = io_reset; // @[:@138799.4 RegFile.scala 76:16:@138806.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@138805.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@138809.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@138803.4]
  assign regs_369_clock = clock; // @[:@138812.4]
  assign regs_369_reset = io_reset; // @[:@138813.4 RegFile.scala 76:16:@138820.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@138819.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@138823.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@138817.4]
  assign regs_370_clock = clock; // @[:@138826.4]
  assign regs_370_reset = io_reset; // @[:@138827.4 RegFile.scala 76:16:@138834.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@138833.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@138837.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@138831.4]
  assign regs_371_clock = clock; // @[:@138840.4]
  assign regs_371_reset = io_reset; // @[:@138841.4 RegFile.scala 76:16:@138848.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@138847.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@138851.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@138845.4]
  assign regs_372_clock = clock; // @[:@138854.4]
  assign regs_372_reset = io_reset; // @[:@138855.4 RegFile.scala 76:16:@138862.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@138861.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@138865.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@138859.4]
  assign regs_373_clock = clock; // @[:@138868.4]
  assign regs_373_reset = io_reset; // @[:@138869.4 RegFile.scala 76:16:@138876.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@138875.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@138879.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@138873.4]
  assign regs_374_clock = clock; // @[:@138882.4]
  assign regs_374_reset = io_reset; // @[:@138883.4 RegFile.scala 76:16:@138890.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@138889.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@138893.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@138887.4]
  assign regs_375_clock = clock; // @[:@138896.4]
  assign regs_375_reset = io_reset; // @[:@138897.4 RegFile.scala 76:16:@138904.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@138903.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@138907.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@138901.4]
  assign regs_376_clock = clock; // @[:@138910.4]
  assign regs_376_reset = io_reset; // @[:@138911.4 RegFile.scala 76:16:@138918.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@138917.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@138921.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@138915.4]
  assign regs_377_clock = clock; // @[:@138924.4]
  assign regs_377_reset = io_reset; // @[:@138925.4 RegFile.scala 76:16:@138932.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@138931.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@138935.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@138929.4]
  assign regs_378_clock = clock; // @[:@138938.4]
  assign regs_378_reset = io_reset; // @[:@138939.4 RegFile.scala 76:16:@138946.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@138945.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@138949.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@138943.4]
  assign regs_379_clock = clock; // @[:@138952.4]
  assign regs_379_reset = io_reset; // @[:@138953.4 RegFile.scala 76:16:@138960.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@138959.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@138963.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@138957.4]
  assign regs_380_clock = clock; // @[:@138966.4]
  assign regs_380_reset = io_reset; // @[:@138967.4 RegFile.scala 76:16:@138974.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@138973.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@138977.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@138971.4]
  assign regs_381_clock = clock; // @[:@138980.4]
  assign regs_381_reset = io_reset; // @[:@138981.4 RegFile.scala 76:16:@138988.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@138987.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@138991.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@138985.4]
  assign regs_382_clock = clock; // @[:@138994.4]
  assign regs_382_reset = io_reset; // @[:@138995.4 RegFile.scala 76:16:@139002.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@139001.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@139005.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@138999.4]
  assign regs_383_clock = clock; // @[:@139008.4]
  assign regs_383_reset = io_reset; // @[:@139009.4 RegFile.scala 76:16:@139016.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@139015.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@139019.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@139013.4]
  assign regs_384_clock = clock; // @[:@139022.4]
  assign regs_384_reset = io_reset; // @[:@139023.4 RegFile.scala 76:16:@139030.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@139029.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@139033.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@139027.4]
  assign regs_385_clock = clock; // @[:@139036.4]
  assign regs_385_reset = io_reset; // @[:@139037.4 RegFile.scala 76:16:@139044.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@139043.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@139047.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@139041.4]
  assign regs_386_clock = clock; // @[:@139050.4]
  assign regs_386_reset = io_reset; // @[:@139051.4 RegFile.scala 76:16:@139058.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@139057.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@139061.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@139055.4]
  assign regs_387_clock = clock; // @[:@139064.4]
  assign regs_387_reset = io_reset; // @[:@139065.4 RegFile.scala 76:16:@139072.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@139071.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@139075.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@139069.4]
  assign regs_388_clock = clock; // @[:@139078.4]
  assign regs_388_reset = io_reset; // @[:@139079.4 RegFile.scala 76:16:@139086.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@139085.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@139089.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@139083.4]
  assign regs_389_clock = clock; // @[:@139092.4]
  assign regs_389_reset = io_reset; // @[:@139093.4 RegFile.scala 76:16:@139100.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@139099.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@139103.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@139097.4]
  assign regs_390_clock = clock; // @[:@139106.4]
  assign regs_390_reset = io_reset; // @[:@139107.4 RegFile.scala 76:16:@139114.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@139113.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@139117.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@139111.4]
  assign regs_391_clock = clock; // @[:@139120.4]
  assign regs_391_reset = io_reset; // @[:@139121.4 RegFile.scala 76:16:@139128.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@139127.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@139131.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@139125.4]
  assign regs_392_clock = clock; // @[:@139134.4]
  assign regs_392_reset = io_reset; // @[:@139135.4 RegFile.scala 76:16:@139142.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@139141.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@139145.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@139139.4]
  assign regs_393_clock = clock; // @[:@139148.4]
  assign regs_393_reset = io_reset; // @[:@139149.4 RegFile.scala 76:16:@139156.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@139155.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@139159.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@139153.4]
  assign regs_394_clock = clock; // @[:@139162.4]
  assign regs_394_reset = io_reset; // @[:@139163.4 RegFile.scala 76:16:@139170.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@139169.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@139173.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@139167.4]
  assign regs_395_clock = clock; // @[:@139176.4]
  assign regs_395_reset = io_reset; // @[:@139177.4 RegFile.scala 76:16:@139184.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@139183.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@139187.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@139181.4]
  assign regs_396_clock = clock; // @[:@139190.4]
  assign regs_396_reset = io_reset; // @[:@139191.4 RegFile.scala 76:16:@139198.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@139197.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@139201.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@139195.4]
  assign regs_397_clock = clock; // @[:@139204.4]
  assign regs_397_reset = io_reset; // @[:@139205.4 RegFile.scala 76:16:@139212.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@139211.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@139215.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@139209.4]
  assign regs_398_clock = clock; // @[:@139218.4]
  assign regs_398_reset = io_reset; // @[:@139219.4 RegFile.scala 76:16:@139226.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@139225.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@139229.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@139223.4]
  assign regs_399_clock = clock; // @[:@139232.4]
  assign regs_399_reset = io_reset; // @[:@139233.4 RegFile.scala 76:16:@139240.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@139239.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@139243.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@139237.4]
  assign regs_400_clock = clock; // @[:@139246.4]
  assign regs_400_reset = io_reset; // @[:@139247.4 RegFile.scala 76:16:@139254.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@139253.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@139257.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@139251.4]
  assign regs_401_clock = clock; // @[:@139260.4]
  assign regs_401_reset = io_reset; // @[:@139261.4 RegFile.scala 76:16:@139268.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@139267.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@139271.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@139265.4]
  assign regs_402_clock = clock; // @[:@139274.4]
  assign regs_402_reset = io_reset; // @[:@139275.4 RegFile.scala 76:16:@139282.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@139281.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@139285.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@139279.4]
  assign regs_403_clock = clock; // @[:@139288.4]
  assign regs_403_reset = io_reset; // @[:@139289.4 RegFile.scala 76:16:@139296.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@139295.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@139299.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@139293.4]
  assign regs_404_clock = clock; // @[:@139302.4]
  assign regs_404_reset = io_reset; // @[:@139303.4 RegFile.scala 76:16:@139310.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@139309.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@139313.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@139307.4]
  assign regs_405_clock = clock; // @[:@139316.4]
  assign regs_405_reset = io_reset; // @[:@139317.4 RegFile.scala 76:16:@139324.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@139323.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@139327.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@139321.4]
  assign regs_406_clock = clock; // @[:@139330.4]
  assign regs_406_reset = io_reset; // @[:@139331.4 RegFile.scala 76:16:@139338.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@139337.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@139341.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@139335.4]
  assign regs_407_clock = clock; // @[:@139344.4]
  assign regs_407_reset = io_reset; // @[:@139345.4 RegFile.scala 76:16:@139352.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@139351.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@139355.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@139349.4]
  assign regs_408_clock = clock; // @[:@139358.4]
  assign regs_408_reset = io_reset; // @[:@139359.4 RegFile.scala 76:16:@139366.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@139365.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@139369.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@139363.4]
  assign regs_409_clock = clock; // @[:@139372.4]
  assign regs_409_reset = io_reset; // @[:@139373.4 RegFile.scala 76:16:@139380.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@139379.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@139383.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@139377.4]
  assign regs_410_clock = clock; // @[:@139386.4]
  assign regs_410_reset = io_reset; // @[:@139387.4 RegFile.scala 76:16:@139394.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@139393.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@139397.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@139391.4]
  assign regs_411_clock = clock; // @[:@139400.4]
  assign regs_411_reset = io_reset; // @[:@139401.4 RegFile.scala 76:16:@139408.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@139407.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@139411.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@139405.4]
  assign regs_412_clock = clock; // @[:@139414.4]
  assign regs_412_reset = io_reset; // @[:@139415.4 RegFile.scala 76:16:@139422.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@139421.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@139425.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@139419.4]
  assign regs_413_clock = clock; // @[:@139428.4]
  assign regs_413_reset = io_reset; // @[:@139429.4 RegFile.scala 76:16:@139436.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@139435.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@139439.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@139433.4]
  assign regs_414_clock = clock; // @[:@139442.4]
  assign regs_414_reset = io_reset; // @[:@139443.4 RegFile.scala 76:16:@139450.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@139449.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@139453.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@139447.4]
  assign regs_415_clock = clock; // @[:@139456.4]
  assign regs_415_reset = io_reset; // @[:@139457.4 RegFile.scala 76:16:@139464.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@139463.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@139467.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@139461.4]
  assign regs_416_clock = clock; // @[:@139470.4]
  assign regs_416_reset = io_reset; // @[:@139471.4 RegFile.scala 76:16:@139478.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@139477.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@139481.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@139475.4]
  assign regs_417_clock = clock; // @[:@139484.4]
  assign regs_417_reset = io_reset; // @[:@139485.4 RegFile.scala 76:16:@139492.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@139491.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@139495.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@139489.4]
  assign regs_418_clock = clock; // @[:@139498.4]
  assign regs_418_reset = io_reset; // @[:@139499.4 RegFile.scala 76:16:@139506.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@139505.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@139509.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@139503.4]
  assign regs_419_clock = clock; // @[:@139512.4]
  assign regs_419_reset = io_reset; // @[:@139513.4 RegFile.scala 76:16:@139520.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@139519.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@139523.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@139517.4]
  assign regs_420_clock = clock; // @[:@139526.4]
  assign regs_420_reset = io_reset; // @[:@139527.4 RegFile.scala 76:16:@139534.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@139533.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@139537.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@139531.4]
  assign regs_421_clock = clock; // @[:@139540.4]
  assign regs_421_reset = io_reset; // @[:@139541.4 RegFile.scala 76:16:@139548.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@139547.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@139551.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@139545.4]
  assign regs_422_clock = clock; // @[:@139554.4]
  assign regs_422_reset = io_reset; // @[:@139555.4 RegFile.scala 76:16:@139562.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@139561.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@139565.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@139559.4]
  assign regs_423_clock = clock; // @[:@139568.4]
  assign regs_423_reset = io_reset; // @[:@139569.4 RegFile.scala 76:16:@139576.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@139575.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@139579.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@139573.4]
  assign regs_424_clock = clock; // @[:@139582.4]
  assign regs_424_reset = io_reset; // @[:@139583.4 RegFile.scala 76:16:@139590.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@139589.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@139593.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@139587.4]
  assign regs_425_clock = clock; // @[:@139596.4]
  assign regs_425_reset = io_reset; // @[:@139597.4 RegFile.scala 76:16:@139604.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@139603.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@139607.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@139601.4]
  assign regs_426_clock = clock; // @[:@139610.4]
  assign regs_426_reset = io_reset; // @[:@139611.4 RegFile.scala 76:16:@139618.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@139617.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@139621.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@139615.4]
  assign regs_427_clock = clock; // @[:@139624.4]
  assign regs_427_reset = io_reset; // @[:@139625.4 RegFile.scala 76:16:@139632.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@139631.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@139635.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@139629.4]
  assign regs_428_clock = clock; // @[:@139638.4]
  assign regs_428_reset = io_reset; // @[:@139639.4 RegFile.scala 76:16:@139646.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@139645.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@139649.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@139643.4]
  assign regs_429_clock = clock; // @[:@139652.4]
  assign regs_429_reset = io_reset; // @[:@139653.4 RegFile.scala 76:16:@139660.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@139659.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@139663.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@139657.4]
  assign regs_430_clock = clock; // @[:@139666.4]
  assign regs_430_reset = io_reset; // @[:@139667.4 RegFile.scala 76:16:@139674.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@139673.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@139677.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@139671.4]
  assign regs_431_clock = clock; // @[:@139680.4]
  assign regs_431_reset = io_reset; // @[:@139681.4 RegFile.scala 76:16:@139688.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@139687.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@139691.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@139685.4]
  assign regs_432_clock = clock; // @[:@139694.4]
  assign regs_432_reset = io_reset; // @[:@139695.4 RegFile.scala 76:16:@139702.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@139701.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@139705.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@139699.4]
  assign regs_433_clock = clock; // @[:@139708.4]
  assign regs_433_reset = io_reset; // @[:@139709.4 RegFile.scala 76:16:@139716.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@139715.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@139719.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@139713.4]
  assign regs_434_clock = clock; // @[:@139722.4]
  assign regs_434_reset = io_reset; // @[:@139723.4 RegFile.scala 76:16:@139730.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@139729.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@139733.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@139727.4]
  assign regs_435_clock = clock; // @[:@139736.4]
  assign regs_435_reset = io_reset; // @[:@139737.4 RegFile.scala 76:16:@139744.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@139743.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@139747.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@139741.4]
  assign regs_436_clock = clock; // @[:@139750.4]
  assign regs_436_reset = io_reset; // @[:@139751.4 RegFile.scala 76:16:@139758.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@139757.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@139761.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@139755.4]
  assign regs_437_clock = clock; // @[:@139764.4]
  assign regs_437_reset = io_reset; // @[:@139765.4 RegFile.scala 76:16:@139772.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@139771.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@139775.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@139769.4]
  assign regs_438_clock = clock; // @[:@139778.4]
  assign regs_438_reset = io_reset; // @[:@139779.4 RegFile.scala 76:16:@139786.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@139785.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@139789.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@139783.4]
  assign regs_439_clock = clock; // @[:@139792.4]
  assign regs_439_reset = io_reset; // @[:@139793.4 RegFile.scala 76:16:@139800.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@139799.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@139803.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@139797.4]
  assign regs_440_clock = clock; // @[:@139806.4]
  assign regs_440_reset = io_reset; // @[:@139807.4 RegFile.scala 76:16:@139814.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@139813.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@139817.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@139811.4]
  assign regs_441_clock = clock; // @[:@139820.4]
  assign regs_441_reset = io_reset; // @[:@139821.4 RegFile.scala 76:16:@139828.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@139827.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@139831.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@139825.4]
  assign regs_442_clock = clock; // @[:@139834.4]
  assign regs_442_reset = io_reset; // @[:@139835.4 RegFile.scala 76:16:@139842.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@139841.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@139845.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@139839.4]
  assign regs_443_clock = clock; // @[:@139848.4]
  assign regs_443_reset = io_reset; // @[:@139849.4 RegFile.scala 76:16:@139856.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@139855.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@139859.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@139853.4]
  assign regs_444_clock = clock; // @[:@139862.4]
  assign regs_444_reset = io_reset; // @[:@139863.4 RegFile.scala 76:16:@139870.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@139869.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@139873.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@139867.4]
  assign regs_445_clock = clock; // @[:@139876.4]
  assign regs_445_reset = io_reset; // @[:@139877.4 RegFile.scala 76:16:@139884.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@139883.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@139887.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@139881.4]
  assign regs_446_clock = clock; // @[:@139890.4]
  assign regs_446_reset = io_reset; // @[:@139891.4 RegFile.scala 76:16:@139898.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@139897.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@139901.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@139895.4]
  assign regs_447_clock = clock; // @[:@139904.4]
  assign regs_447_reset = io_reset; // @[:@139905.4 RegFile.scala 76:16:@139912.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@139911.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@139915.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@139909.4]
  assign regs_448_clock = clock; // @[:@139918.4]
  assign regs_448_reset = io_reset; // @[:@139919.4 RegFile.scala 76:16:@139926.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@139925.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@139929.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@139923.4]
  assign regs_449_clock = clock; // @[:@139932.4]
  assign regs_449_reset = io_reset; // @[:@139933.4 RegFile.scala 76:16:@139940.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@139939.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@139943.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@139937.4]
  assign regs_450_clock = clock; // @[:@139946.4]
  assign regs_450_reset = io_reset; // @[:@139947.4 RegFile.scala 76:16:@139954.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@139953.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@139957.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@139951.4]
  assign regs_451_clock = clock; // @[:@139960.4]
  assign regs_451_reset = io_reset; // @[:@139961.4 RegFile.scala 76:16:@139968.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@139967.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@139971.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@139965.4]
  assign regs_452_clock = clock; // @[:@139974.4]
  assign regs_452_reset = io_reset; // @[:@139975.4 RegFile.scala 76:16:@139982.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@139981.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@139985.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@139979.4]
  assign regs_453_clock = clock; // @[:@139988.4]
  assign regs_453_reset = io_reset; // @[:@139989.4 RegFile.scala 76:16:@139996.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@139995.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@139999.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@139993.4]
  assign regs_454_clock = clock; // @[:@140002.4]
  assign regs_454_reset = io_reset; // @[:@140003.4 RegFile.scala 76:16:@140010.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@140009.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@140013.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@140007.4]
  assign regs_455_clock = clock; // @[:@140016.4]
  assign regs_455_reset = io_reset; // @[:@140017.4 RegFile.scala 76:16:@140024.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@140023.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@140027.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@140021.4]
  assign regs_456_clock = clock; // @[:@140030.4]
  assign regs_456_reset = io_reset; // @[:@140031.4 RegFile.scala 76:16:@140038.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@140037.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@140041.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@140035.4]
  assign regs_457_clock = clock; // @[:@140044.4]
  assign regs_457_reset = io_reset; // @[:@140045.4 RegFile.scala 76:16:@140052.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@140051.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@140055.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@140049.4]
  assign regs_458_clock = clock; // @[:@140058.4]
  assign regs_458_reset = io_reset; // @[:@140059.4 RegFile.scala 76:16:@140066.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@140065.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@140069.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@140063.4]
  assign regs_459_clock = clock; // @[:@140072.4]
  assign regs_459_reset = io_reset; // @[:@140073.4 RegFile.scala 76:16:@140080.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@140079.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@140083.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@140077.4]
  assign regs_460_clock = clock; // @[:@140086.4]
  assign regs_460_reset = io_reset; // @[:@140087.4 RegFile.scala 76:16:@140094.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@140093.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@140097.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@140091.4]
  assign regs_461_clock = clock; // @[:@140100.4]
  assign regs_461_reset = io_reset; // @[:@140101.4 RegFile.scala 76:16:@140108.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@140107.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@140111.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@140105.4]
  assign regs_462_clock = clock; // @[:@140114.4]
  assign regs_462_reset = io_reset; // @[:@140115.4 RegFile.scala 76:16:@140122.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@140121.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@140125.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@140119.4]
  assign regs_463_clock = clock; // @[:@140128.4]
  assign regs_463_reset = io_reset; // @[:@140129.4 RegFile.scala 76:16:@140136.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@140135.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@140139.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@140133.4]
  assign regs_464_clock = clock; // @[:@140142.4]
  assign regs_464_reset = io_reset; // @[:@140143.4 RegFile.scala 76:16:@140150.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@140149.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@140153.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@140147.4]
  assign regs_465_clock = clock; // @[:@140156.4]
  assign regs_465_reset = io_reset; // @[:@140157.4 RegFile.scala 76:16:@140164.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@140163.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@140167.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@140161.4]
  assign regs_466_clock = clock; // @[:@140170.4]
  assign regs_466_reset = io_reset; // @[:@140171.4 RegFile.scala 76:16:@140178.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@140177.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@140181.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@140175.4]
  assign regs_467_clock = clock; // @[:@140184.4]
  assign regs_467_reset = io_reset; // @[:@140185.4 RegFile.scala 76:16:@140192.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@140191.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@140195.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@140189.4]
  assign regs_468_clock = clock; // @[:@140198.4]
  assign regs_468_reset = io_reset; // @[:@140199.4 RegFile.scala 76:16:@140206.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@140205.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@140209.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@140203.4]
  assign regs_469_clock = clock; // @[:@140212.4]
  assign regs_469_reset = io_reset; // @[:@140213.4 RegFile.scala 76:16:@140220.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@140219.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@140223.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@140217.4]
  assign regs_470_clock = clock; // @[:@140226.4]
  assign regs_470_reset = io_reset; // @[:@140227.4 RegFile.scala 76:16:@140234.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@140233.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@140237.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@140231.4]
  assign regs_471_clock = clock; // @[:@140240.4]
  assign regs_471_reset = io_reset; // @[:@140241.4 RegFile.scala 76:16:@140248.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@140247.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@140251.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@140245.4]
  assign regs_472_clock = clock; // @[:@140254.4]
  assign regs_472_reset = io_reset; // @[:@140255.4 RegFile.scala 76:16:@140262.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@140261.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@140265.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@140259.4]
  assign regs_473_clock = clock; // @[:@140268.4]
  assign regs_473_reset = io_reset; // @[:@140269.4 RegFile.scala 76:16:@140276.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@140275.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@140279.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@140273.4]
  assign regs_474_clock = clock; // @[:@140282.4]
  assign regs_474_reset = io_reset; // @[:@140283.4 RegFile.scala 76:16:@140290.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@140289.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@140293.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@140287.4]
  assign regs_475_clock = clock; // @[:@140296.4]
  assign regs_475_reset = io_reset; // @[:@140297.4 RegFile.scala 76:16:@140304.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@140303.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@140307.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@140301.4]
  assign regs_476_clock = clock; // @[:@140310.4]
  assign regs_476_reset = io_reset; // @[:@140311.4 RegFile.scala 76:16:@140318.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@140317.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@140321.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@140315.4]
  assign regs_477_clock = clock; // @[:@140324.4]
  assign regs_477_reset = io_reset; // @[:@140325.4 RegFile.scala 76:16:@140332.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@140331.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@140335.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@140329.4]
  assign regs_478_clock = clock; // @[:@140338.4]
  assign regs_478_reset = io_reset; // @[:@140339.4 RegFile.scala 76:16:@140346.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@140345.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@140349.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@140343.4]
  assign regs_479_clock = clock; // @[:@140352.4]
  assign regs_479_reset = io_reset; // @[:@140353.4 RegFile.scala 76:16:@140360.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@140359.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@140363.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@140357.4]
  assign regs_480_clock = clock; // @[:@140366.4]
  assign regs_480_reset = io_reset; // @[:@140367.4 RegFile.scala 76:16:@140374.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@140373.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@140377.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@140371.4]
  assign regs_481_clock = clock; // @[:@140380.4]
  assign regs_481_reset = io_reset; // @[:@140381.4 RegFile.scala 76:16:@140388.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@140387.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@140391.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@140385.4]
  assign regs_482_clock = clock; // @[:@140394.4]
  assign regs_482_reset = io_reset; // @[:@140395.4 RegFile.scala 76:16:@140402.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@140401.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@140405.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@140399.4]
  assign regs_483_clock = clock; // @[:@140408.4]
  assign regs_483_reset = io_reset; // @[:@140409.4 RegFile.scala 76:16:@140416.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@140415.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@140419.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@140413.4]
  assign regs_484_clock = clock; // @[:@140422.4]
  assign regs_484_reset = io_reset; // @[:@140423.4 RegFile.scala 76:16:@140430.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@140429.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@140433.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@140427.4]
  assign regs_485_clock = clock; // @[:@140436.4]
  assign regs_485_reset = io_reset; // @[:@140437.4 RegFile.scala 76:16:@140444.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@140443.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@140447.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@140441.4]
  assign regs_486_clock = clock; // @[:@140450.4]
  assign regs_486_reset = io_reset; // @[:@140451.4 RegFile.scala 76:16:@140458.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@140457.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@140461.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@140455.4]
  assign regs_487_clock = clock; // @[:@140464.4]
  assign regs_487_reset = io_reset; // @[:@140465.4 RegFile.scala 76:16:@140472.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@140471.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@140475.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@140469.4]
  assign regs_488_clock = clock; // @[:@140478.4]
  assign regs_488_reset = io_reset; // @[:@140479.4 RegFile.scala 76:16:@140486.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@140485.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@140489.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@140483.4]
  assign regs_489_clock = clock; // @[:@140492.4]
  assign regs_489_reset = io_reset; // @[:@140493.4 RegFile.scala 76:16:@140500.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@140499.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@140503.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@140497.4]
  assign regs_490_clock = clock; // @[:@140506.4]
  assign regs_490_reset = io_reset; // @[:@140507.4 RegFile.scala 76:16:@140514.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@140513.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@140517.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@140511.4]
  assign regs_491_clock = clock; // @[:@140520.4]
  assign regs_491_reset = io_reset; // @[:@140521.4 RegFile.scala 76:16:@140528.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@140527.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@140531.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@140525.4]
  assign regs_492_clock = clock; // @[:@140534.4]
  assign regs_492_reset = io_reset; // @[:@140535.4 RegFile.scala 76:16:@140542.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@140541.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@140545.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@140539.4]
  assign regs_493_clock = clock; // @[:@140548.4]
  assign regs_493_reset = io_reset; // @[:@140549.4 RegFile.scala 76:16:@140556.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@140555.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@140559.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@140553.4]
  assign regs_494_clock = clock; // @[:@140562.4]
  assign regs_494_reset = io_reset; // @[:@140563.4 RegFile.scala 76:16:@140570.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@140569.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@140573.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@140567.4]
  assign regs_495_clock = clock; // @[:@140576.4]
  assign regs_495_reset = io_reset; // @[:@140577.4 RegFile.scala 76:16:@140584.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@140583.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@140587.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@140581.4]
  assign regs_496_clock = clock; // @[:@140590.4]
  assign regs_496_reset = io_reset; // @[:@140591.4 RegFile.scala 76:16:@140598.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@140597.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@140601.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@140595.4]
  assign regs_497_clock = clock; // @[:@140604.4]
  assign regs_497_reset = io_reset; // @[:@140605.4 RegFile.scala 76:16:@140612.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@140611.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@140615.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@140609.4]
  assign regs_498_clock = clock; // @[:@140618.4]
  assign regs_498_reset = io_reset; // @[:@140619.4 RegFile.scala 76:16:@140626.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@140625.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@140629.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@140623.4]
  assign regs_499_clock = clock; // @[:@140632.4]
  assign regs_499_reset = io_reset; // @[:@140633.4 RegFile.scala 76:16:@140640.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@140639.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@140643.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@140637.4]
  assign regs_500_clock = clock; // @[:@140646.4]
  assign regs_500_reset = io_reset; // @[:@140647.4 RegFile.scala 76:16:@140654.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@140653.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@140657.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@140651.4]
  assign regs_501_clock = clock; // @[:@140660.4]
  assign regs_501_reset = io_reset; // @[:@140661.4 RegFile.scala 76:16:@140668.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@140667.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@140671.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@140665.4]
  assign regs_502_clock = clock; // @[:@140674.4]
  assign regs_502_reset = io_reset; // @[:@140675.4 RegFile.scala 76:16:@140682.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@140681.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@140685.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@140679.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@141194.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@141195.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@141196.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@141197.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@141198.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@141199.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@141200.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@141201.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@141202.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@141203.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@141204.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@141205.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@141206.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@141207.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@141208.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@141209.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@141210.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@141211.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@141212.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@141213.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@141214.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@141215.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@141216.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@141217.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@141218.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@141219.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@141220.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@141221.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@141222.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@141223.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@141224.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@141225.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@141226.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@141227.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@141228.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@141229.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@141230.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@141231.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@141232.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@141233.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@141234.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@141235.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@141236.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@141237.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@141238.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@141239.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@141240.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@141241.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@141242.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@141243.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@141244.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@141245.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@141246.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@141247.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@141248.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@141249.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@141250.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@141251.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@141252.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@141253.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@141254.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@141255.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@141256.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@141257.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@141258.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@141259.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@141260.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@141261.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@141262.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@141263.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@141264.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@141265.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@141266.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@141267.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@141268.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@141269.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@141270.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@141271.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@141272.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@141273.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@141274.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@141275.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@141276.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@141277.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@141278.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@141279.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@141280.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@141281.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@141282.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@141283.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@141284.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@141285.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@141286.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@141287.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@141288.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@141289.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@141290.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@141291.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@141292.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@141293.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@141294.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@141295.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@141296.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@141297.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@141298.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@141299.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@141300.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@141301.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@141302.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@141303.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@141304.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@141305.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@141306.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@141307.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@141308.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@141309.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@141310.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@141311.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@141312.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@141313.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@141314.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@141315.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@141316.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@141317.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@141318.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@141319.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@141320.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@141321.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@141322.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@141323.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@141324.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@141325.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@141326.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@141327.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@141328.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@141329.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@141330.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@141331.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@141332.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@141333.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@141334.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@141335.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@141336.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@141337.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@141338.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@141339.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@141340.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@141341.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@141342.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@141343.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@141344.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@141345.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@141346.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@141347.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@141348.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@141349.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@141350.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@141351.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@141352.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@141353.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@141354.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@141355.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@141356.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@141357.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@141358.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@141359.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@141360.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@141361.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@141362.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@141363.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@141364.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@141365.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@141366.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@141367.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@141368.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@141369.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@141370.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@141371.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@141372.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@141373.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@141374.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@141375.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@141376.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@141377.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@141378.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@141379.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@141380.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@141381.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@141382.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@141383.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@141384.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@141385.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@141386.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@141387.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@141388.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@141389.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@141390.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@141391.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@141392.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@141393.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@141394.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@141395.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@141396.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@141397.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@141398.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@141399.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@141400.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@141401.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@141402.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@141403.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@141404.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@141405.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@141406.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@141407.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@141408.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@141409.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@141410.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@141411.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@141412.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@141413.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@141414.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@141415.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@141416.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@141417.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@141418.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@141419.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@141420.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@141421.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@141422.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@141423.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@141424.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@141425.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@141426.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@141427.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@141428.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@141429.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@141430.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@141431.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@141432.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@141433.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@141434.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@141435.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@141436.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@141437.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@141438.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@141439.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@141440.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@141441.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@141442.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@141443.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@141444.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@141445.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@141446.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@141447.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@141448.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@141449.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@141450.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@141451.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@141452.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@141453.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@141454.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@141455.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@141456.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@141457.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@141458.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@141459.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@141460.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@141461.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@141462.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@141463.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@141464.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@141465.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@141466.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@141467.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@141468.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@141469.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@141470.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@141471.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@141472.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@141473.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@141474.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@141475.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@141476.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@141477.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@141478.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@141479.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@141480.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@141481.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@141482.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@141483.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@141484.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@141485.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@141486.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@141487.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@141488.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@141489.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@141490.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@141491.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@141492.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@141493.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@141494.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@141495.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@141496.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@141497.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@141498.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@141499.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@141500.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@141501.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@141502.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@141503.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@141504.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@141505.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@141506.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@141507.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@141508.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@141509.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@141510.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@141511.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@141512.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@141513.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@141514.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@141515.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@141516.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@141517.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@141518.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@141519.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@141520.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@141521.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@141522.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@141523.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@141524.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@141525.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@141526.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@141527.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@141528.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@141529.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@141530.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@141531.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@141532.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@141533.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@141534.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@141535.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@141536.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@141537.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@141538.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@141539.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@141540.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@141541.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@141542.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@141543.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@141544.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@141545.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@141546.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@141547.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@141548.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@141549.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@141550.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@141551.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@141552.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@141553.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@141554.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@141555.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@141556.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@141557.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@141558.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@141559.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@141560.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@141561.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@141562.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@141563.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@141564.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@141565.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@141566.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@141567.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@141568.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@141569.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@141570.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@141571.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@141572.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@141573.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@141574.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@141575.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@141576.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@141577.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@141578.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@141579.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@141580.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@141581.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@141582.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@141583.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@141584.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@141585.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@141586.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@141587.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@141588.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@141589.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@141590.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@141591.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@141592.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@141593.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@141594.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@141595.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@141596.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@141597.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@141598.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@141599.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@141600.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@141601.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@141602.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@141603.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@141604.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@141605.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@141606.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@141607.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@141608.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@141609.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@141610.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@141611.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@141612.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@141613.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@141614.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@141615.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@141616.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@141617.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@141618.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@141619.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@141620.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@141621.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@141622.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@141623.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@141624.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@141625.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@141626.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@141627.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@141628.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@141629.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@141630.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@141631.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@141632.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@141633.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@141634.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@141635.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@141636.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@141637.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@141638.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@141639.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@141640.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@141641.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@141642.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@141643.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@141644.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@141645.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@141646.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@141647.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@141648.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@141649.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@141650.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@141651.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@141652.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@141653.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@141654.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@141655.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@141656.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@141657.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@141658.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@141659.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@141660.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@141661.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@141662.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@141663.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@141664.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@141665.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@141666.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@141667.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@141668.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@141669.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@141670.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@141671.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@141672.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@141673.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@141674.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@141675.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@141676.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@141677.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@141678.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@141679.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@141680.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@141681.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@141682.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@141683.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@141684.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@141685.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@141686.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@141687.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@141688.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@141689.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@141690.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@141691.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@141692.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@141693.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@141694.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@141695.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@141696.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@141697.4]
endmodule
module RetimeWrapper_923( // @[:@141721.2]
  input         clock, // @[:@141722.4]
  input         reset, // @[:@141723.4]
  input  [39:0] io_in, // @[:@141724.4]
  output [39:0] io_out // @[:@141724.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@141726.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@141726.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@141726.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@141726.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@141726.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@141726.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@141726.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@141739.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@141738.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@141737.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@141736.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@141735.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@141733.4]
endmodule
module FringeFF_503( // @[:@141741.2]
  input         clock, // @[:@141742.4]
  input         reset, // @[:@141743.4]
  input  [39:0] io_in, // @[:@141744.4]
  output [39:0] io_out, // @[:@141744.4]
  input         io_enable // @[:@141744.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@141747.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@141747.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@141747.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@141747.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@141752.4 package.scala 96:25:@141753.4]
  RetimeWrapper_923 RetimeWrapper ( // @[package.scala 93:22:@141747.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@141752.4 package.scala 96:25:@141753.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@141764.4]
  assign RetimeWrapper_clock = clock; // @[:@141748.4]
  assign RetimeWrapper_reset = reset; // @[:@141749.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@141750.4]
endmodule
module FringeCounter( // @[:@141766.2]
  input   clock, // @[:@141767.4]
  input   reset, // @[:@141768.4]
  input   io_enable, // @[:@141769.4]
  output  io_done // @[:@141769.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@141771.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@141771.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@141771.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@141771.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@141771.4]
  wire [40:0] count; // @[Cat.scala 30:58:@141778.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@141779.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@141780.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@141781.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@141783.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@141771.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@141778.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@141779.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@141780.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@141781.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@141783.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@141794.4]
  assign reg$_clock = clock; // @[:@141772.4]
  assign reg$_reset = reset; // @[:@141773.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@141785.6 FringeCounter.scala 37:15:@141788.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@141776.4]
endmodule
module FringeFF_504( // @[:@141828.2]
  input   clock, // @[:@141829.4]
  input   reset, // @[:@141830.4]
  input   io_in, // @[:@141831.4]
  input   io_reset, // @[:@141831.4]
  output  io_out, // @[:@141831.4]
  input   io_enable // @[:@141831.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@141834.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@141834.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@141834.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@141834.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@141834.4]
  wire  _T_18; // @[package.scala 96:25:@141839.4 package.scala 96:25:@141840.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@141845.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@141834.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@141839.4 package.scala 96:25:@141840.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@141845.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@141851.4]
  assign RetimeWrapper_clock = clock; // @[:@141835.4]
  assign RetimeWrapper_reset = reset; // @[:@141836.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@141838.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@141837.4]
endmodule
module Depulser( // @[:@141853.2]
  input   clock, // @[:@141854.4]
  input   reset, // @[:@141855.4]
  input   io_in, // @[:@141856.4]
  input   io_rst, // @[:@141856.4]
  output  io_out // @[:@141856.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@141858.4]
  wire  r_reset; // @[Depulser.scala 14:17:@141858.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@141858.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@141858.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@141858.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@141858.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@141858.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@141867.4]
  assign r_clock = clock; // @[:@141859.4]
  assign r_reset = reset; // @[:@141860.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@141862.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@141866.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@141865.4]
endmodule
module Fringe( // @[:@141869.2]
  input         clock, // @[:@141870.4]
  input         reset, // @[:@141871.4]
  input  [31:0] io_raddr, // @[:@141872.4]
  input         io_wen, // @[:@141872.4]
  input  [31:0] io_waddr, // @[:@141872.4]
  input  [63:0] io_wdata, // @[:@141872.4]
  output [63:0] io_rdata, // @[:@141872.4]
  output        io_enable, // @[:@141872.4]
  input         io_done, // @[:@141872.4]
  output        io_reset, // @[:@141872.4]
  output [63:0] io_argIns_0, // @[:@141872.4]
  output [63:0] io_argIns_1, // @[:@141872.4]
  input         io_argOuts_0_valid, // @[:@141872.4]
  input  [63:0] io_argOuts_0_bits, // @[:@141872.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@141872.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@141872.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@141872.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@141872.4]
  output        io_memStreams_stores_0_data_ready, // @[:@141872.4]
  input         io_memStreams_stores_0_data_valid, // @[:@141872.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@141872.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@141872.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@141872.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@141872.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@141872.4]
  input         io_dram_0_cmd_ready, // @[:@141872.4]
  output        io_dram_0_cmd_valid, // @[:@141872.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@141872.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@141872.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@141872.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@141872.4]
  input         io_dram_0_wdata_ready, // @[:@141872.4]
  output        io_dram_0_wdata_valid, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@141872.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@141872.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@141872.4]
  output        io_dram_0_rresp_ready, // @[:@141872.4]
  output        io_dram_0_wresp_ready, // @[:@141872.4]
  input         io_dram_0_wresp_valid, // @[:@141872.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@141872.4]
  input         io_dram_1_cmd_ready, // @[:@141872.4]
  output        io_dram_1_cmd_valid, // @[:@141872.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@141872.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@141872.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@141872.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@141872.4]
  input         io_dram_1_wdata_ready, // @[:@141872.4]
  output        io_dram_1_wdata_valid, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@141872.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@141872.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@141872.4]
  output        io_dram_1_rresp_ready, // @[:@141872.4]
  output        io_dram_1_wresp_ready, // @[:@141872.4]
  input         io_dram_1_wresp_valid, // @[:@141872.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@141872.4]
  input         io_dram_2_cmd_ready, // @[:@141872.4]
  output        io_dram_2_cmd_valid, // @[:@141872.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@141872.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@141872.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@141872.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@141872.4]
  input         io_dram_2_wdata_ready, // @[:@141872.4]
  output        io_dram_2_wdata_valid, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@141872.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@141872.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@141872.4]
  output        io_dram_2_rresp_ready, // @[:@141872.4]
  output        io_dram_2_wresp_ready, // @[:@141872.4]
  input         io_dram_2_wresp_valid, // @[:@141872.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@141872.4]
  input         io_dram_3_cmd_ready, // @[:@141872.4]
  output        io_dram_3_cmd_valid, // @[:@141872.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@141872.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@141872.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@141872.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@141872.4]
  input         io_dram_3_wdata_ready, // @[:@141872.4]
  output        io_dram_3_wdata_valid, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@141872.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@141872.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@141872.4]
  output        io_dram_3_rresp_ready, // @[:@141872.4]
  output        io_dram_3_wresp_ready, // @[:@141872.4]
  input         io_dram_3_wresp_valid, // @[:@141872.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@141872.4]
  input         io_heap_0_req_valid, // @[:@141872.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@141872.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@141872.4]
  output        io_heap_0_resp_valid, // @[:@141872.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@141872.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@141872.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@141878.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@141878.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@141878.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@141878.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@142871.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@142871.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@142871.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@143831.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@143831.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@143831.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@144791.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@144791.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@144791.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@144791.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@145751.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@145751.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@145751.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@145751.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@145751.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@145751.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@145751.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@145751.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@145751.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@145751.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@145751.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@145751.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@145760.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@145760.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@145760.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@145760.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@145760.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@145760.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@145760.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@145760.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@145760.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@147810.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@147810.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@147810.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@147810.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@147829.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@147829.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@147829.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@147829.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@147829.4]
  wire [63:0] _T_1020; // @[:@147787.4 :@147788.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@147789.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@147791.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@147793.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@147795.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@147797.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@147799.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@147801.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@147837.4]
  reg  _T_1047; // @[package.scala 152:20:@147840.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@147842.4]
  wire  _T_1049; // @[package.scala 153:8:@147843.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@147847.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@147848.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@147851.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@147852.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@147854.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@147855.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@147857.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@147860.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@147839.4 Fringe.scala 163:24:@147858.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@147839.4 Fringe.scala 162:28:@147856.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@147861.4]
  wire  alloc; // @[Fringe.scala 202:38:@149491.4]
  wire  dealloc; // @[Fringe.scala 203:40:@149492.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@149493.4]
  reg  _T_1572; // @[package.scala 152:20:@149494.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@149496.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@141878.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@142871.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@143831.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@144791.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@145751.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@145760.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@147810.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@147829.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@147787.4 :@147788.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@147789.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@147791.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@147793.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@147795.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@147797.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@147799.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@147801.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@147837.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@147842.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@147843.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@147847.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@147848.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@147851.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@147852.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@147854.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@147855.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@147857.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@147860.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@147839.4 Fringe.scala 163:24:@147858.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@147839.4 Fringe.scala 162:28:@147856.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@147861.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@149491.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@149492.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@149493.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@149496.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@147785.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@147805.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@147806.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@147827.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@147828.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@142797.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@142793.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@142788.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@142787.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@148989.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@148988.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@148987.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@148985.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@148984.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@148982.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@148966.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@148967.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@148968.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@148969.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@148970.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@148971.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@148972.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@148973.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@148974.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@148975.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@148976.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@148977.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@148978.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@148979.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@148980.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@148981.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@148902.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@148903.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@148904.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@148905.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@148906.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@148907.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@148908.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@148909.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@148910.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@148911.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@148912.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@148913.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@148914.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@148915.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@148916.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@148917.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@148918.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@148919.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@148920.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@148921.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@148922.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@148923.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@148924.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@148925.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@148926.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@148927.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@148928.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@148929.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@148930.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@148931.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@148932.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@148933.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@148934.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@148935.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@148936.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@148937.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@148938.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@148939.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@148940.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@148941.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@148942.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@148943.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@148944.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@148945.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@148946.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@148947.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@148948.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@148949.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@148950.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@148951.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@148952.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@148953.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@148954.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@148955.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@148956.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@148957.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@148958.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@148959.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@148960.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@148961.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@148962.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@148963.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@148964.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@148965.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@148901.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@148900.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@148881.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@149101.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@149100.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@149099.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@149097.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@149096.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@149094.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@149078.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@149079.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@149080.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@149081.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@149082.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@149083.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@149084.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@149085.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@149086.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@149087.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@149088.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@149089.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@149090.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@149091.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@149092.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@149093.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@149014.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@149015.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@149016.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@149017.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@149018.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@149019.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@149020.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@149021.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@149022.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@149023.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@149024.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@149025.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@149026.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@149027.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@149028.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@149029.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@149030.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@149031.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@149032.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@149033.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@149034.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@149035.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@149036.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@149037.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@149038.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@149039.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@149040.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@149041.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@149042.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@149043.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@149044.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@149045.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@149046.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@149047.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@149048.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@149049.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@149050.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@149051.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@149052.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@149053.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@149054.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@149055.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@149056.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@149057.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@149058.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@149059.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@149060.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@149061.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@149062.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@149063.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@149064.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@149065.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@149066.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@149067.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@149068.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@149069.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@149070.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@149071.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@149072.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@149073.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@149074.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@149075.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@149076.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@149077.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@149013.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@149012.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@148993.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@149213.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@149212.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@149211.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@149209.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@149208.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@149206.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@149190.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@149191.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@149192.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@149193.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@149194.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@149195.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@149196.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@149197.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@149198.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@149199.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@149200.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@149201.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@149202.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@149203.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@149204.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@149205.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@149126.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@149127.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@149128.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@149129.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@149130.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@149131.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@149132.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@149133.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@149134.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@149135.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@149136.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@149137.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@149138.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@149139.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@149140.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@149141.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@149142.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@149143.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@149144.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@149145.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@149146.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@149147.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@149148.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@149149.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@149150.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@149151.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@149152.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@149153.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@149154.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@149155.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@149156.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@149157.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@149158.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@149159.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@149160.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@149161.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@149162.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@149163.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@149164.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@149165.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@149166.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@149167.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@149168.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@149169.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@149170.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@149171.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@149172.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@149173.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@149174.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@149175.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@149176.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@149177.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@149178.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@149179.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@149180.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@149181.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@149182.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@149183.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@149184.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@149185.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@149186.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@149187.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@149188.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@149189.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@149125.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@149124.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@149105.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@149325.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@149324.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@149323.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@149321.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@149320.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@149318.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@149302.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@149303.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@149304.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@149305.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@149306.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@149307.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@149308.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@149309.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@149310.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@149311.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@149312.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@149313.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@149314.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@149315.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@149316.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@149317.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@149238.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@149239.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@149240.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@149241.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@149242.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@149243.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@149244.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@149245.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@149246.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@149247.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@149248.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@149249.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@149250.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@149251.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@149252.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@149253.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@149254.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@149255.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@149256.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@149257.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@149258.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@149259.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@149260.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@149261.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@149262.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@149263.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@149264.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@149265.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@149266.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@149267.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@149268.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@149269.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@149270.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@149271.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@149272.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@149273.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@149274.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@149275.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@149276.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@149277.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@149278.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@149279.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@149280.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@149281.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@149282.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@149283.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@149284.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@149285.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@149286.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@149287.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@149288.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@149289.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@149290.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@149291.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@149292.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@149293.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@149294.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@149295.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@149296.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@149297.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@149298.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@149299.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@149300.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@149301.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@149237.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@149236.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@149217.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@145756.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@145755.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@145754.4]
  assign dramArbs_0_clock = clock; // @[:@141879.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@141880.4 Fringe.scala 187:30:@148871.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148875.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@142796.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@142795.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@142794.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@142792.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@142791.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@142790.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@142789.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@148990.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@148983.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@148880.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@148879.4]
  assign dramArbs_1_clock = clock; // @[:@142872.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@142873.4 Fringe.scala 187:30:@148872.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148876.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@149102.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@149095.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@148992.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@148991.4]
  assign dramArbs_2_clock = clock; // @[:@143832.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@143833.4 Fringe.scala 187:30:@148873.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148877.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@149214.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@149207.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@149104.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@149103.4]
  assign dramArbs_3_clock = clock; // @[:@144792.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@144793.4 Fringe.scala 187:30:@148874.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148878.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@149326.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@149319.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@149216.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@149215.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@145759.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@145758.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@145757.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@149498.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@149499.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@149500.4]
  assign regs_clock = clock; // @[:@145761.4]
  assign regs_reset = reset; // @[:@145762.4 Fringe.scala 139:14:@147809.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@147781.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@147783.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@147782.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@147784.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@147807.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@147859.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@147863.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@147866.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@147865.4]
  assign timeoutCtr_clock = clock; // @[:@147811.4]
  assign timeoutCtr_reset = reset; // @[:@147812.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@147826.4]
  assign depulser_clock = clock; // @[:@147830.4]
  assign depulser_reset = reset; // @[:@147831.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@147836.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@147838.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@149515.2]
  input         clock, // @[:@149516.4]
  input         reset, // @[:@149517.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@149518.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@149518.4]
  input         io_S_AXI_AWVALID, // @[:@149518.4]
  output        io_S_AXI_AWREADY, // @[:@149518.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@149518.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@149518.4]
  input         io_S_AXI_ARVALID, // @[:@149518.4]
  output        io_S_AXI_ARREADY, // @[:@149518.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@149518.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@149518.4]
  input         io_S_AXI_WVALID, // @[:@149518.4]
  output        io_S_AXI_WREADY, // @[:@149518.4]
  output [31:0] io_S_AXI_RDATA, // @[:@149518.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@149518.4]
  output        io_S_AXI_RVALID, // @[:@149518.4]
  input         io_S_AXI_RREADY, // @[:@149518.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@149518.4]
  output        io_S_AXI_BVALID, // @[:@149518.4]
  input         io_S_AXI_BREADY, // @[:@149518.4]
  output [31:0] io_raddr, // @[:@149518.4]
  output        io_wen, // @[:@149518.4]
  output [31:0] io_waddr, // @[:@149518.4]
  output [31:0] io_wdata, // @[:@149518.4]
  input  [31:0] io_rdata // @[:@149518.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@149520.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149544.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149540.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149536.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@149535.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@149534.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149533.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@149531.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149530.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@149552.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@149555.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@149553.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@149554.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@149556.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@149551.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@149548.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@149547.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@149546.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149545.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@149543.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@149542.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149541.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@149539.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@149538.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149537.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149532.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149529.4]
endmodule
module MAGToAXI4Bridge( // @[:@149558.2]
  output         io_in_cmd_ready, // @[:@149561.4]
  input          io_in_cmd_valid, // @[:@149561.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@149561.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@149561.4]
  input          io_in_cmd_bits_isWr, // @[:@149561.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@149561.4]
  output         io_in_wdata_ready, // @[:@149561.4]
  input          io_in_wdata_valid, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@149561.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@149561.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@149561.4]
  input          io_in_wdata_bits_wlast, // @[:@149561.4]
  input          io_in_rresp_ready, // @[:@149561.4]
  input          io_in_wresp_ready, // @[:@149561.4]
  output         io_in_wresp_valid, // @[:@149561.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@149561.4]
  output [31:0]  io_M_AXI_AWID, // @[:@149561.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@149561.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@149561.4]
  output         io_M_AXI_AWVALID, // @[:@149561.4]
  input          io_M_AXI_AWREADY, // @[:@149561.4]
  output [31:0]  io_M_AXI_ARID, // @[:@149561.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@149561.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@149561.4]
  output         io_M_AXI_ARVALID, // @[:@149561.4]
  input          io_M_AXI_ARREADY, // @[:@149561.4]
  output [511:0] io_M_AXI_WDATA, // @[:@149561.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@149561.4]
  output         io_M_AXI_WLAST, // @[:@149561.4]
  output         io_M_AXI_WVALID, // @[:@149561.4]
  input          io_M_AXI_WREADY, // @[:@149561.4]
  output         io_M_AXI_RREADY, // @[:@149561.4]
  input  [31:0]  io_M_AXI_BID, // @[:@149561.4]
  input          io_M_AXI_BVALID, // @[:@149561.4]
  output         io_M_AXI_BREADY // @[:@149561.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@149718.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@149719.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@149720.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@149728.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@149755.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@149760.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@149771.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@149780.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@149789.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@149798.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@149807.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@149816.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@149824.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@149718.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@149719.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@149720.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@149728.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@149755.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@149760.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@149771.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@149780.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@149789.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@149798.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@149807.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@149816.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@149824.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@149732.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@149829.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@149882.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@149884.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@149733.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@149734.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@149738.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@149746.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@149716.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@149717.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@149721.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@149730.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@149762.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@149826.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@149827.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@149828.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@149879.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@149880.4]
endmodule
module FringeZynq( // @[:@150870.2]
  input          clock, // @[:@150871.4]
  input          reset, // @[:@150872.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@150873.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@150873.4]
  input          io_S_AXI_AWVALID, // @[:@150873.4]
  output         io_S_AXI_AWREADY, // @[:@150873.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@150873.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@150873.4]
  input          io_S_AXI_ARVALID, // @[:@150873.4]
  output         io_S_AXI_ARREADY, // @[:@150873.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@150873.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@150873.4]
  input          io_S_AXI_WVALID, // @[:@150873.4]
  output         io_S_AXI_WREADY, // @[:@150873.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@150873.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@150873.4]
  output         io_S_AXI_RVALID, // @[:@150873.4]
  input          io_S_AXI_RREADY, // @[:@150873.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@150873.4]
  output         io_S_AXI_BVALID, // @[:@150873.4]
  input          io_S_AXI_BREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@150873.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@150873.4]
  output         io_M_AXI_0_AWVALID, // @[:@150873.4]
  input          io_M_AXI_0_AWREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@150873.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@150873.4]
  output         io_M_AXI_0_ARVALID, // @[:@150873.4]
  input          io_M_AXI_0_ARREADY, // @[:@150873.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@150873.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@150873.4]
  output         io_M_AXI_0_WLAST, // @[:@150873.4]
  output         io_M_AXI_0_WVALID, // @[:@150873.4]
  input          io_M_AXI_0_WREADY, // @[:@150873.4]
  output         io_M_AXI_0_RREADY, // @[:@150873.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@150873.4]
  input          io_M_AXI_0_BVALID, // @[:@150873.4]
  output         io_M_AXI_0_BREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@150873.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@150873.4]
  output         io_M_AXI_1_AWVALID, // @[:@150873.4]
  input          io_M_AXI_1_AWREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@150873.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@150873.4]
  output         io_M_AXI_1_ARVALID, // @[:@150873.4]
  input          io_M_AXI_1_ARREADY, // @[:@150873.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@150873.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@150873.4]
  output         io_M_AXI_1_WLAST, // @[:@150873.4]
  output         io_M_AXI_1_WVALID, // @[:@150873.4]
  input          io_M_AXI_1_WREADY, // @[:@150873.4]
  output         io_M_AXI_1_RREADY, // @[:@150873.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@150873.4]
  input          io_M_AXI_1_BVALID, // @[:@150873.4]
  output         io_M_AXI_1_BREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@150873.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@150873.4]
  output         io_M_AXI_2_AWVALID, // @[:@150873.4]
  input          io_M_AXI_2_AWREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@150873.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@150873.4]
  output         io_M_AXI_2_ARVALID, // @[:@150873.4]
  input          io_M_AXI_2_ARREADY, // @[:@150873.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@150873.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@150873.4]
  output         io_M_AXI_2_WLAST, // @[:@150873.4]
  output         io_M_AXI_2_WVALID, // @[:@150873.4]
  input          io_M_AXI_2_WREADY, // @[:@150873.4]
  output         io_M_AXI_2_RREADY, // @[:@150873.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@150873.4]
  input          io_M_AXI_2_BVALID, // @[:@150873.4]
  output         io_M_AXI_2_BREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@150873.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@150873.4]
  output         io_M_AXI_3_AWVALID, // @[:@150873.4]
  input          io_M_AXI_3_AWREADY, // @[:@150873.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@150873.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@150873.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@150873.4]
  output         io_M_AXI_3_ARVALID, // @[:@150873.4]
  input          io_M_AXI_3_ARREADY, // @[:@150873.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@150873.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@150873.4]
  output         io_M_AXI_3_WLAST, // @[:@150873.4]
  output         io_M_AXI_3_WVALID, // @[:@150873.4]
  input          io_M_AXI_3_WREADY, // @[:@150873.4]
  output         io_M_AXI_3_RREADY, // @[:@150873.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@150873.4]
  input          io_M_AXI_3_BVALID, // @[:@150873.4]
  output         io_M_AXI_3_BREADY, // @[:@150873.4]
  output         io_enable, // @[:@150873.4]
  input          io_done, // @[:@150873.4]
  output         io_reset, // @[:@150873.4]
  output [63:0]  io_argIns_0, // @[:@150873.4]
  output [63:0]  io_argIns_1, // @[:@150873.4]
  input          io_argOuts_0_valid, // @[:@150873.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@150873.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@150873.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@150873.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@150873.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@150873.4]
  output         io_memStreams_stores_0_data_ready, // @[:@150873.4]
  input          io_memStreams_stores_0_data_valid, // @[:@150873.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@150873.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@150873.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@150873.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@150873.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@150873.4]
  input          io_heap_0_req_valid, // @[:@150873.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@150873.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@150873.4]
  output         io_heap_0_resp_valid, // @[:@150873.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@150873.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@150873.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@151344.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@151344.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@151344.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@152250.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@152250.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@152250.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@152250.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@152250.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@152250.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@152250.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@152250.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152400.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152400.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152400.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152400.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152400.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152400.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152400.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152556.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152556.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152556.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152556.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152556.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152556.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152556.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152712.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152712.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152712.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152712.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152712.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152712.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152712.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152868.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152868.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152868.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152868.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152868.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152868.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152868.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152868.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@151344.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@152250.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@152400.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@152556.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@152712.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@152868.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@152268.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@152264.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@152260.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@152259.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@152258.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@152257.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@152255.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@152254.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@152555.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@152553.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@152552.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@152545.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@152543.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@152541.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@152540.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@152533.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152531.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152530.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152529.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152528.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152520.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152515.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@152711.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@152709.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@152708.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@152701.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@152699.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@152697.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@152696.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@152689.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152687.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152686.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152685.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152684.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152676.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152671.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@152867.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@152865.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@152864.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@152857.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@152855.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@152853.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@152852.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@152845.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152843.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152842.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152841.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152840.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152832.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152827.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@153023.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@153021.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@153020.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@153013.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@153011.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@153009.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@153008.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@153001.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152999.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152998.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152997.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152996.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152988.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152983.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@152278.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@152282.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@152283.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@152284.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@152371.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@152367.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@152362.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@152361.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@152396.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@152395.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@152394.4]
  assign fringeCommon_clock = clock; // @[:@151345.4]
  assign fringeCommon_reset = reset; // @[:@151346.4 FringeZynq.scala 117:22:@152281.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@152272.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@152273.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@152274.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@152275.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@152279.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@152286.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@152285.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@152370.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@152369.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@152368.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@152366.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@152365.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@152364.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@152363.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152514.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152507.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152404.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152403.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152670.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152663.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152560.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152559.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152826.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152819.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152716.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152715.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152982.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152975.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152872.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152871.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@152399.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@152398.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@152397.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@152251.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@152252.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@152271.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@152270.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@152269.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@152267.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@152266.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@152265.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@152263.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@152262.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@152261.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@152256.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@152253.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@152276.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@152513.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152512.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@152511.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152509.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152508.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@152506.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152490.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152491.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152492.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152493.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152494.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152495.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152496.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152497.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152498.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152499.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152500.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152501.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152502.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152503.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152504.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152505.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152426.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152427.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152428.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152429.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152430.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152431.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152432.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152433.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152434.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152435.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152436.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152437.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152438.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152439.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152440.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152441.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152442.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152443.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152444.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152445.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152446.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152447.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152448.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152449.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152450.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152451.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152452.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152453.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152454.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152455.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152456.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152457.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152458.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152459.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152460.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152461.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152462.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152463.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152464.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152465.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152466.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152467.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152468.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152469.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152470.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152471.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152472.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152473.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152474.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152475.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152476.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152477.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152478.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152479.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152480.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152481.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152482.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152483.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152484.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152485.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152486.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152487.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152488.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152489.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152425.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@152424.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@152405.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@152544.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@152532.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@152527.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@152519.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@152516.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@152669.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152668.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@152667.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152665.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152664.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@152662.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152646.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152647.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152648.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152649.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152650.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152651.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152652.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152653.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152654.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152655.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152656.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152657.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152658.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152659.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152660.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152661.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152582.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152583.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152584.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152585.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152586.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152587.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152588.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152589.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152590.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152591.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152592.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152593.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152594.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152595.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152596.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152597.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152598.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152599.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152600.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152601.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152602.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152603.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152604.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152605.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152606.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152607.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152608.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152609.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152610.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152611.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152612.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152613.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152614.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152615.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152616.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152617.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152618.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152619.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152620.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152621.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152622.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152623.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152624.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152625.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152626.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152627.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152628.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152629.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152630.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152631.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152632.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152633.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152634.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152635.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152636.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152637.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152638.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152639.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152640.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152641.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152642.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152643.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152644.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152645.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152581.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@152580.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@152561.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@152700.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@152688.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@152683.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@152675.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@152672.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@152825.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152824.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@152823.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152821.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152820.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@152818.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152802.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152803.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152804.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152805.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152806.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152807.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152808.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152809.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152810.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152811.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152812.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152813.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152814.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152815.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152816.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152817.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152738.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152739.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152740.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152741.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152742.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152743.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152744.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152745.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152746.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152747.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152748.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152749.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152750.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152751.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152752.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152753.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152754.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152755.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152756.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152757.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152758.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152759.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152760.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152761.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152762.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152763.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152764.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152765.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152766.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152767.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152768.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152769.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152770.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152771.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152772.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152773.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152774.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152775.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152776.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152777.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152778.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152779.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152780.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152781.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152782.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152783.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152784.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152785.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152786.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152787.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152788.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152789.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152790.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152791.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152792.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152793.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152794.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152795.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152796.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152797.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152798.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152799.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152800.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152801.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152737.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@152736.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@152717.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@152856.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@152844.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@152839.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@152831.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@152828.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@152981.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152980.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@152979.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152977.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152976.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@152974.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152958.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152959.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152960.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152961.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152962.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152963.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152964.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152965.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152966.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152967.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152968.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152969.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152970.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152971.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152972.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152973.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152894.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152895.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152896.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152897.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152898.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152899.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152900.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152901.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152902.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152903.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152904.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152905.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152906.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152907.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152908.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152909.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152910.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152911.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152912.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152913.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152914.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152915.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152916.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152917.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152918.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152919.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152920.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152921.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152922.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152923.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152924.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152925.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152926.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152927.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152928.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152929.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152930.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152931.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152932.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152933.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152934.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152935.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152936.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152937.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152938.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152939.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152940.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152941.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152942.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152943.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152944.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152945.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152946.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152947.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152948.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152949.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152950.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152951.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152952.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152953.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152954.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152955.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152956.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152957.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152893.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@152892.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@152873.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@153012.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@153000.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@152995.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@152987.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@152984.4]
endmodule
module SpatialIP( // @[:@153025.2]
  input          clock, // @[:@153026.4]
  input          reset, // @[:@153027.4]
  input          io_raddr, // @[:@153028.4]
  input          io_wen, // @[:@153028.4]
  input          io_waddr, // @[:@153028.4]
  input          io_wdata, // @[:@153028.4]
  output         io_rdata, // @[:@153028.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@153028.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@153028.4]
  input          io_S_AXI_AWVALID, // @[:@153028.4]
  output         io_S_AXI_AWREADY, // @[:@153028.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@153028.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@153028.4]
  input          io_S_AXI_ARVALID, // @[:@153028.4]
  output         io_S_AXI_ARREADY, // @[:@153028.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@153028.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@153028.4]
  input          io_S_AXI_WVALID, // @[:@153028.4]
  output         io_S_AXI_WREADY, // @[:@153028.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@153028.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@153028.4]
  output         io_S_AXI_RVALID, // @[:@153028.4]
  input          io_S_AXI_RREADY, // @[:@153028.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@153028.4]
  output         io_S_AXI_BVALID, // @[:@153028.4]
  input          io_S_AXI_BREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@153028.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@153028.4]
  output         io_M_AXI_0_AWLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@153028.4]
  output         io_M_AXI_0_AWVALID, // @[:@153028.4]
  input          io_M_AXI_0_AWREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@153028.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@153028.4]
  output         io_M_AXI_0_ARLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@153028.4]
  output         io_M_AXI_0_ARVALID, // @[:@153028.4]
  input          io_M_AXI_0_ARREADY, // @[:@153028.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@153028.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@153028.4]
  output         io_M_AXI_0_WLAST, // @[:@153028.4]
  output         io_M_AXI_0_WVALID, // @[:@153028.4]
  input          io_M_AXI_0_WREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@153028.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@153028.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@153028.4]
  input          io_M_AXI_0_RLAST, // @[:@153028.4]
  input          io_M_AXI_0_RVALID, // @[:@153028.4]
  output         io_M_AXI_0_RREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@153028.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@153028.4]
  input          io_M_AXI_0_BVALID, // @[:@153028.4]
  output         io_M_AXI_0_BREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@153028.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@153028.4]
  output         io_M_AXI_1_AWLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@153028.4]
  output         io_M_AXI_1_AWVALID, // @[:@153028.4]
  input          io_M_AXI_1_AWREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@153028.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@153028.4]
  output         io_M_AXI_1_ARLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@153028.4]
  output         io_M_AXI_1_ARVALID, // @[:@153028.4]
  input          io_M_AXI_1_ARREADY, // @[:@153028.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@153028.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@153028.4]
  output         io_M_AXI_1_WLAST, // @[:@153028.4]
  output         io_M_AXI_1_WVALID, // @[:@153028.4]
  input          io_M_AXI_1_WREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@153028.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@153028.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@153028.4]
  input          io_M_AXI_1_RLAST, // @[:@153028.4]
  input          io_M_AXI_1_RVALID, // @[:@153028.4]
  output         io_M_AXI_1_RREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@153028.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@153028.4]
  input          io_M_AXI_1_BVALID, // @[:@153028.4]
  output         io_M_AXI_1_BREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@153028.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@153028.4]
  output         io_M_AXI_2_AWLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@153028.4]
  output         io_M_AXI_2_AWVALID, // @[:@153028.4]
  input          io_M_AXI_2_AWREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@153028.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@153028.4]
  output         io_M_AXI_2_ARLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@153028.4]
  output         io_M_AXI_2_ARVALID, // @[:@153028.4]
  input          io_M_AXI_2_ARREADY, // @[:@153028.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@153028.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@153028.4]
  output         io_M_AXI_2_WLAST, // @[:@153028.4]
  output         io_M_AXI_2_WVALID, // @[:@153028.4]
  input          io_M_AXI_2_WREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@153028.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@153028.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@153028.4]
  input          io_M_AXI_2_RLAST, // @[:@153028.4]
  input          io_M_AXI_2_RVALID, // @[:@153028.4]
  output         io_M_AXI_2_RREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@153028.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@153028.4]
  input          io_M_AXI_2_BVALID, // @[:@153028.4]
  output         io_M_AXI_2_BREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@153028.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@153028.4]
  output         io_M_AXI_3_AWLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@153028.4]
  output         io_M_AXI_3_AWVALID, // @[:@153028.4]
  input          io_M_AXI_3_AWREADY, // @[:@153028.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@153028.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@153028.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@153028.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@153028.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@153028.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@153028.4]
  output         io_M_AXI_3_ARLOCK, // @[:@153028.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@153028.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@153028.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@153028.4]
  output         io_M_AXI_3_ARVALID, // @[:@153028.4]
  input          io_M_AXI_3_ARREADY, // @[:@153028.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@153028.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@153028.4]
  output         io_M_AXI_3_WLAST, // @[:@153028.4]
  output         io_M_AXI_3_WVALID, // @[:@153028.4]
  input          io_M_AXI_3_WREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@153028.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@153028.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@153028.4]
  input          io_M_AXI_3_RLAST, // @[:@153028.4]
  input          io_M_AXI_3_RVALID, // @[:@153028.4]
  output         io_M_AXI_3_RREADY, // @[:@153028.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@153028.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@153028.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@153028.4]
  input          io_M_AXI_3_BVALID, // @[:@153028.4]
  output         io_M_AXI_3_BREADY, // @[:@153028.4]
  input          io_TOP_AXI_AWID, // @[:@153028.4]
  input          io_TOP_AXI_AWUSER, // @[:@153028.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@153028.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@153028.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@153028.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@153028.4]
  input          io_TOP_AXI_AWLOCK, // @[:@153028.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@153028.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@153028.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@153028.4]
  input          io_TOP_AXI_AWVALID, // @[:@153028.4]
  input          io_TOP_AXI_AWREADY, // @[:@153028.4]
  input          io_TOP_AXI_ARID, // @[:@153028.4]
  input          io_TOP_AXI_ARUSER, // @[:@153028.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@153028.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@153028.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@153028.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@153028.4]
  input          io_TOP_AXI_ARLOCK, // @[:@153028.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@153028.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@153028.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@153028.4]
  input          io_TOP_AXI_ARVALID, // @[:@153028.4]
  input          io_TOP_AXI_ARREADY, // @[:@153028.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@153028.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@153028.4]
  input          io_TOP_AXI_WLAST, // @[:@153028.4]
  input          io_TOP_AXI_WVALID, // @[:@153028.4]
  input          io_TOP_AXI_WREADY, // @[:@153028.4]
  input          io_TOP_AXI_RID, // @[:@153028.4]
  input          io_TOP_AXI_RUSER, // @[:@153028.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@153028.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@153028.4]
  input          io_TOP_AXI_RLAST, // @[:@153028.4]
  input          io_TOP_AXI_RVALID, // @[:@153028.4]
  input          io_TOP_AXI_RREADY, // @[:@153028.4]
  input          io_TOP_AXI_BID, // @[:@153028.4]
  input          io_TOP_AXI_BUSER, // @[:@153028.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@153028.4]
  input          io_TOP_AXI_BVALID, // @[:@153028.4]
  input          io_TOP_AXI_BREADY, // @[:@153028.4]
  input          io_DWIDTH_AXI_AWID, // @[:@153028.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@153028.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@153028.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@153028.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@153028.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@153028.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@153028.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@153028.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@153028.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@153028.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@153028.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@153028.4]
  input          io_DWIDTH_AXI_ARID, // @[:@153028.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@153028.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@153028.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@153028.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@153028.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@153028.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@153028.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@153028.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@153028.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@153028.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@153028.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@153028.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@153028.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@153028.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@153028.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@153028.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@153028.4]
  input          io_DWIDTH_AXI_RID, // @[:@153028.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@153028.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@153028.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@153028.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@153028.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@153028.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@153028.4]
  input          io_DWIDTH_AXI_BID, // @[:@153028.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@153028.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@153028.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@153028.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@153028.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@153028.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@153028.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@153028.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@153028.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@153028.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@153028.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@153028.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@153028.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@153028.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@153028.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@153028.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@153028.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@153028.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@153028.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@153028.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@153028.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@153028.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@153028.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@153028.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@153028.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@153028.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@153028.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@153028.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@153028.4]
  input          io_PROTOCOL_AXI_RID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@153028.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@153028.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@153028.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@153028.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@153028.4]
  input          io_PROTOCOL_AXI_BID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@153028.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@153028.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@153028.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@153028.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@153028.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@153028.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@153028.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@153028.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@153028.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@153028.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@153028.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@153028.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@153028.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@153028.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@153028.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@153028.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@153028.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@153028.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@153028.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@153028.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@153028.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@153028.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@153028.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@153028.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@153030.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@153030.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@153030.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@153030.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@153030.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@153030.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@153030.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@153030.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@153030.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@153030.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@153172.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@153172.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@153172.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@153172.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@153172.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@153172.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@153172.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@153030.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@153172.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@153190.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@153186.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@153182.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@153181.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@153180.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@153179.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@153177.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@153176.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@153234.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153233.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@153232.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@153231.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153230.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153229.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153228.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153227.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153226.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153225.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@153224.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@153222.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153221.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@153220.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@153219.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153218.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153217.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153216.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153215.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153214.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153213.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@153212.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@153210.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@153209.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@153208.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@153207.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@153199.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@153194.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@153275.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153274.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@153273.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@153272.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153271.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153270.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153269.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153268.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153267.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153266.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@153265.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@153263.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153262.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@153261.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@153260.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153259.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153258.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153257.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153256.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153255.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153254.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@153253.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@153251.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@153250.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@153249.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@153248.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@153240.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@153235.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@153316.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153315.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@153314.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@153313.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153312.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153311.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153310.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153309.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153308.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153307.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@153306.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@153304.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153303.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@153302.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@153301.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153300.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153299.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153298.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153297.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153296.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153295.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@153294.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@153292.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@153291.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@153290.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@153289.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@153281.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@153276.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@153357.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153356.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@153355.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@153354.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153353.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153352.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153351.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153350.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153349.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153348.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@153347.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@153345.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153344.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@153343.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@153342.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153341.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153340.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153339.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153338.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153337.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153336.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@153335.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@153333.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@153332.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@153331.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@153330.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@153322.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@153317.4]
  assign accel_clock = clock; // @[:@153031.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@153032.4 Zynq.scala 54:17:@153646.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@153641.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@153634.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@153629.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@153613.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@153614.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@153615.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@153616.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@153617.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@153618.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@153619.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@153620.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@153621.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@153622.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@153623.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@153624.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@153625.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@153626.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@153627.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@153628.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@153612.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@153608.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@153603.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@153602.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@153601.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@153582.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@153566.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@153567.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@153568.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@153569.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@153570.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@153571.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@153572.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@153573.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@153574.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@153575.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@153576.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@153577.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@153578.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@153579.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@153580.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@153581.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@153565.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@153530.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@153529.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@153637.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@153636.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@153635.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@153523.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@153524.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@153527.4]
  assign FringeZynq_clock = clock; // @[:@153173.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@153174.4 Zynq.scala 53:18:@153645.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@153193.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@153192.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@153191.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@153189.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@153188.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@153187.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@153185.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@153184.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@153183.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@153178.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@153175.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@153223.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@153211.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@153206.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@153198.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@153195.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@153264.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@153252.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@153247.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@153239.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@153236.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@153305.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@153293.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@153288.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@153280.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@153277.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@153346.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@153334.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@153329.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@153321.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@153318.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@153642.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@153526.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@153525.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@153611.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@153610.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@153609.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@153607.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@153606.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@153605.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@153604.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@153640.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@153639.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@153638.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




