module FIFO(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  input  [15:0] I_8,
  input  [15:0] I_9,
  input  [15:0] I_10,
  input  [15:0] I_11,
  input  [15:0] I_12,
  input  [15:0] I_13,
  input  [15:0] I_14,
  input  [15:0] I_15,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7,
  output [15:0] O_8,
  output [15:0] O_9,
  output [15:0] O_10,
  output [15:0] O_11,
  output [15:0] O_12,
  output [15:0] O_13,
  output [15:0] O_14,
  output [15:0] O_15
);
  reg [15:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [15:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [15:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [15:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [15:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [15:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [15:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [15:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [15:0] _T__8; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [15:0] _T__9; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [15:0] _T__10; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [15:0] _T__11; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [15:0] _T__12; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [15:0] _T__13; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [15:0] _T__14; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [15:0] _T__15; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_16;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
  assign O_8 = _T__8; // @[FIFO.scala 14:7]
  assign O_9 = _T__9; // @[FIFO.scala 14:7]
  assign O_10 = _T__10; // @[FIFO.scala 14:7]
  assign O_11 = _T__11; // @[FIFO.scala 14:7]
  assign O_12 = _T__12; // @[FIFO.scala 14:7]
  assign O_13 = _T__13; // @[FIFO.scala 14:7]
  assign O_14 = _T__14; // @[FIFO.scala 14:7]
  assign O_15 = _T__15; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__9 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__10 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__11 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__12 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__13 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__14 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__15 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    _T__8 <= I_8;
    _T__9 <= I_9;
    _T__10 <= I_10;
    _T__11 <= I_11;
    _T__12 <= I_12;
    _T__13 <= I_13;
    _T__14 <= I_14;
    _T__15 <= I_15;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input         clock,
  input         RE,
  input  [6:0]  RADDR,
  output [15:0] RDATA,
  input         WE,
  input  [6:0]  WADDR,
  input  [15:0] WDATA
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [15:0] ram [0:119]; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_0;
  wire [15:0] ram__T_8_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram__T_8_addr; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_1;
  wire [15:0] ram__T_2_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram__T_2_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_8_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [6:0] ram__T_8_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [6:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [7:0] _T; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_126; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_127; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_128; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_129; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_130; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_131; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_132; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_133; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_134; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_135; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_136; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_137; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_138; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_139; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_140; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_141; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_142; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_143; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_144; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_145; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_146; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_147; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_148; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_149; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_150; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_151; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_152; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_153; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_154; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_155; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_156; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_157; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_158; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_159; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_160; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_161; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_162; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_163; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_164; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_165; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_166; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_167; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_168; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_169; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_170; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_171; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_172; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_173; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_174; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_175; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_176; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_177; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_178; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_179; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_180; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_181; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_182; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_183; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_184; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_185; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_186; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_187; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_188; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_189; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_190; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_191; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_192; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_193; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_194; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_195; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_196; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_197; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_198; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_199; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_200; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_201; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_202; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_203; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_204; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_205; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_206; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_207; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_208; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_209; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_210; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_211; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_212; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_213; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_214; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_215; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_216; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_217; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_218; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_219; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_220; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_221; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_222; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_223; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_224; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_225; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_226; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_227; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_228; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_229; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_230; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_231; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_232; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_233; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_234; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_235; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_236; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_237; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_238; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_239; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_240; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_241; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_242; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_243; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_244; // @[RAM_ST.scala 32:46]
  wire [7:0] _T_3; // @[RAM_ST.scala 32:46]
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_8_addr = ram__T_8_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_8_data = ram[ram__T_8_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_8_data = ram__T_8_addr >= 7'h78 ? _RAND_1[15:0] : ram[ram__T_8_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_2_data = WDATA;
  assign ram__T_2_addr = _T[6:0];
  assign ram__T_2_mask = 1'h1;
  assign ram__T_2_en = write_elem_counter_valid;
  assign _GEN_1 = 7'h1 == WADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 7'h2 == WADDR ? 7'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 7'h3 == WADDR ? 7'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 7'h4 == WADDR ? 7'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 7'h5 == WADDR ? 7'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 7'h6 == WADDR ? 7'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 7'h7 == WADDR ? 7'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 7'h8 == WADDR ? 7'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 7'h9 == WADDR ? 7'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 7'ha == WADDR ? 7'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 7'hb == WADDR ? 7'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 7'hc == WADDR ? 7'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 7'hd == WADDR ? 7'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 7'he == WADDR ? 7'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 7'hf == WADDR ? 7'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 7'h10 == WADDR ? 7'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 7'h11 == WADDR ? 7'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 7'h12 == WADDR ? 7'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 7'h13 == WADDR ? 7'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 7'h14 == WADDR ? 7'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 7'h15 == WADDR ? 7'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 7'h16 == WADDR ? 7'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 7'h17 == WADDR ? 7'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 7'h18 == WADDR ? 7'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 7'h19 == WADDR ? 7'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 7'h1a == WADDR ? 7'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 7'h1b == WADDR ? 7'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 7'h1c == WADDR ? 7'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 7'h1d == WADDR ? 7'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 7'h1e == WADDR ? 7'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 7'h1f == WADDR ? 7'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 7'h20 == WADDR ? 7'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 7'h21 == WADDR ? 7'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 7'h22 == WADDR ? 7'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 7'h23 == WADDR ? 7'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 7'h24 == WADDR ? 7'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 7'h25 == WADDR ? 7'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 7'h26 == WADDR ? 7'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 7'h27 == WADDR ? 7'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 7'h28 == WADDR ? 7'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 7'h29 == WADDR ? 7'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 7'h2a == WADDR ? 7'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 7'h2b == WADDR ? 7'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 7'h2c == WADDR ? 7'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 7'h2d == WADDR ? 7'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 7'h2e == WADDR ? 7'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 7'h2f == WADDR ? 7'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 7'h30 == WADDR ? 7'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 7'h31 == WADDR ? 7'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 7'h32 == WADDR ? 7'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 7'h33 == WADDR ? 7'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 7'h34 == WADDR ? 7'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 7'h35 == WADDR ? 7'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 7'h36 == WADDR ? 7'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 7'h37 == WADDR ? 7'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 7'h38 == WADDR ? 7'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 7'h39 == WADDR ? 7'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 7'h3a == WADDR ? 7'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 7'h3b == WADDR ? 7'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 7'h3c == WADDR ? 7'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 7'h3d == WADDR ? 7'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 7'h3e == WADDR ? 7'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 7'h3f == WADDR ? 7'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 7'h40 == WADDR ? 7'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 7'h41 == WADDR ? 7'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 7'h42 == WADDR ? 7'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 7'h43 == WADDR ? 7'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 7'h44 == WADDR ? 7'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 7'h45 == WADDR ? 7'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 7'h46 == WADDR ? 7'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 7'h47 == WADDR ? 7'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 7'h48 == WADDR ? 7'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 7'h49 == WADDR ? 7'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 7'h4a == WADDR ? 7'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 7'h4b == WADDR ? 7'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 7'h4c == WADDR ? 7'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 7'h4d == WADDR ? 7'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 7'h4e == WADDR ? 7'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 7'h4f == WADDR ? 7'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 7'h50 == WADDR ? 7'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 7'h51 == WADDR ? 7'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 7'h52 == WADDR ? 7'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 7'h53 == WADDR ? 7'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 7'h54 == WADDR ? 7'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 7'h55 == WADDR ? 7'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 7'h56 == WADDR ? 7'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 7'h57 == WADDR ? 7'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 7'h58 == WADDR ? 7'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 7'h59 == WADDR ? 7'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 7'h5a == WADDR ? 7'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 7'h5b == WADDR ? 7'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 7'h5c == WADDR ? 7'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 7'h5d == WADDR ? 7'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 7'h5e == WADDR ? 7'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 7'h5f == WADDR ? 7'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 7'h60 == WADDR ? 7'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 7'h61 == WADDR ? 7'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 7'h62 == WADDR ? 7'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 7'h63 == WADDR ? 7'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 7'h64 == WADDR ? 7'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 7'h65 == WADDR ? 7'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 7'h66 == WADDR ? 7'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 7'h67 == WADDR ? 7'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 7'h68 == WADDR ? 7'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 7'h69 == WADDR ? 7'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 7'h6a == WADDR ? 7'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 7'h6b == WADDR ? 7'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 7'h6c == WADDR ? 7'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 7'h6d == WADDR ? 7'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 7'h6e == WADDR ? 7'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 7'h6f == WADDR ? 7'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 7'h70 == WADDR ? 7'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 7'h71 == WADDR ? 7'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 7'h72 == WADDR ? 7'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 7'h73 == WADDR ? 7'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 7'h74 == WADDR ? 7'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 7'h75 == WADDR ? 7'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 7'h76 == WADDR ? 7'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 7'h77 == WADDR ? 7'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_119}; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 7'h1 == RADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_127 = 7'h2 == RADDR ? 7'h2 : _GEN_126; // @[RAM_ST.scala 32:46]
  assign _GEN_128 = 7'h3 == RADDR ? 7'h3 : _GEN_127; // @[RAM_ST.scala 32:46]
  assign _GEN_129 = 7'h4 == RADDR ? 7'h4 : _GEN_128; // @[RAM_ST.scala 32:46]
  assign _GEN_130 = 7'h5 == RADDR ? 7'h5 : _GEN_129; // @[RAM_ST.scala 32:46]
  assign _GEN_131 = 7'h6 == RADDR ? 7'h6 : _GEN_130; // @[RAM_ST.scala 32:46]
  assign _GEN_132 = 7'h7 == RADDR ? 7'h7 : _GEN_131; // @[RAM_ST.scala 32:46]
  assign _GEN_133 = 7'h8 == RADDR ? 7'h8 : _GEN_132; // @[RAM_ST.scala 32:46]
  assign _GEN_134 = 7'h9 == RADDR ? 7'h9 : _GEN_133; // @[RAM_ST.scala 32:46]
  assign _GEN_135 = 7'ha == RADDR ? 7'ha : _GEN_134; // @[RAM_ST.scala 32:46]
  assign _GEN_136 = 7'hb == RADDR ? 7'hb : _GEN_135; // @[RAM_ST.scala 32:46]
  assign _GEN_137 = 7'hc == RADDR ? 7'hc : _GEN_136; // @[RAM_ST.scala 32:46]
  assign _GEN_138 = 7'hd == RADDR ? 7'hd : _GEN_137; // @[RAM_ST.scala 32:46]
  assign _GEN_139 = 7'he == RADDR ? 7'he : _GEN_138; // @[RAM_ST.scala 32:46]
  assign _GEN_140 = 7'hf == RADDR ? 7'hf : _GEN_139; // @[RAM_ST.scala 32:46]
  assign _GEN_141 = 7'h10 == RADDR ? 7'h10 : _GEN_140; // @[RAM_ST.scala 32:46]
  assign _GEN_142 = 7'h11 == RADDR ? 7'h11 : _GEN_141; // @[RAM_ST.scala 32:46]
  assign _GEN_143 = 7'h12 == RADDR ? 7'h12 : _GEN_142; // @[RAM_ST.scala 32:46]
  assign _GEN_144 = 7'h13 == RADDR ? 7'h13 : _GEN_143; // @[RAM_ST.scala 32:46]
  assign _GEN_145 = 7'h14 == RADDR ? 7'h14 : _GEN_144; // @[RAM_ST.scala 32:46]
  assign _GEN_146 = 7'h15 == RADDR ? 7'h15 : _GEN_145; // @[RAM_ST.scala 32:46]
  assign _GEN_147 = 7'h16 == RADDR ? 7'h16 : _GEN_146; // @[RAM_ST.scala 32:46]
  assign _GEN_148 = 7'h17 == RADDR ? 7'h17 : _GEN_147; // @[RAM_ST.scala 32:46]
  assign _GEN_149 = 7'h18 == RADDR ? 7'h18 : _GEN_148; // @[RAM_ST.scala 32:46]
  assign _GEN_150 = 7'h19 == RADDR ? 7'h19 : _GEN_149; // @[RAM_ST.scala 32:46]
  assign _GEN_151 = 7'h1a == RADDR ? 7'h1a : _GEN_150; // @[RAM_ST.scala 32:46]
  assign _GEN_152 = 7'h1b == RADDR ? 7'h1b : _GEN_151; // @[RAM_ST.scala 32:46]
  assign _GEN_153 = 7'h1c == RADDR ? 7'h1c : _GEN_152; // @[RAM_ST.scala 32:46]
  assign _GEN_154 = 7'h1d == RADDR ? 7'h1d : _GEN_153; // @[RAM_ST.scala 32:46]
  assign _GEN_155 = 7'h1e == RADDR ? 7'h1e : _GEN_154; // @[RAM_ST.scala 32:46]
  assign _GEN_156 = 7'h1f == RADDR ? 7'h1f : _GEN_155; // @[RAM_ST.scala 32:46]
  assign _GEN_157 = 7'h20 == RADDR ? 7'h20 : _GEN_156; // @[RAM_ST.scala 32:46]
  assign _GEN_158 = 7'h21 == RADDR ? 7'h21 : _GEN_157; // @[RAM_ST.scala 32:46]
  assign _GEN_159 = 7'h22 == RADDR ? 7'h22 : _GEN_158; // @[RAM_ST.scala 32:46]
  assign _GEN_160 = 7'h23 == RADDR ? 7'h23 : _GEN_159; // @[RAM_ST.scala 32:46]
  assign _GEN_161 = 7'h24 == RADDR ? 7'h24 : _GEN_160; // @[RAM_ST.scala 32:46]
  assign _GEN_162 = 7'h25 == RADDR ? 7'h25 : _GEN_161; // @[RAM_ST.scala 32:46]
  assign _GEN_163 = 7'h26 == RADDR ? 7'h26 : _GEN_162; // @[RAM_ST.scala 32:46]
  assign _GEN_164 = 7'h27 == RADDR ? 7'h27 : _GEN_163; // @[RAM_ST.scala 32:46]
  assign _GEN_165 = 7'h28 == RADDR ? 7'h28 : _GEN_164; // @[RAM_ST.scala 32:46]
  assign _GEN_166 = 7'h29 == RADDR ? 7'h29 : _GEN_165; // @[RAM_ST.scala 32:46]
  assign _GEN_167 = 7'h2a == RADDR ? 7'h2a : _GEN_166; // @[RAM_ST.scala 32:46]
  assign _GEN_168 = 7'h2b == RADDR ? 7'h2b : _GEN_167; // @[RAM_ST.scala 32:46]
  assign _GEN_169 = 7'h2c == RADDR ? 7'h2c : _GEN_168; // @[RAM_ST.scala 32:46]
  assign _GEN_170 = 7'h2d == RADDR ? 7'h2d : _GEN_169; // @[RAM_ST.scala 32:46]
  assign _GEN_171 = 7'h2e == RADDR ? 7'h2e : _GEN_170; // @[RAM_ST.scala 32:46]
  assign _GEN_172 = 7'h2f == RADDR ? 7'h2f : _GEN_171; // @[RAM_ST.scala 32:46]
  assign _GEN_173 = 7'h30 == RADDR ? 7'h30 : _GEN_172; // @[RAM_ST.scala 32:46]
  assign _GEN_174 = 7'h31 == RADDR ? 7'h31 : _GEN_173; // @[RAM_ST.scala 32:46]
  assign _GEN_175 = 7'h32 == RADDR ? 7'h32 : _GEN_174; // @[RAM_ST.scala 32:46]
  assign _GEN_176 = 7'h33 == RADDR ? 7'h33 : _GEN_175; // @[RAM_ST.scala 32:46]
  assign _GEN_177 = 7'h34 == RADDR ? 7'h34 : _GEN_176; // @[RAM_ST.scala 32:46]
  assign _GEN_178 = 7'h35 == RADDR ? 7'h35 : _GEN_177; // @[RAM_ST.scala 32:46]
  assign _GEN_179 = 7'h36 == RADDR ? 7'h36 : _GEN_178; // @[RAM_ST.scala 32:46]
  assign _GEN_180 = 7'h37 == RADDR ? 7'h37 : _GEN_179; // @[RAM_ST.scala 32:46]
  assign _GEN_181 = 7'h38 == RADDR ? 7'h38 : _GEN_180; // @[RAM_ST.scala 32:46]
  assign _GEN_182 = 7'h39 == RADDR ? 7'h39 : _GEN_181; // @[RAM_ST.scala 32:46]
  assign _GEN_183 = 7'h3a == RADDR ? 7'h3a : _GEN_182; // @[RAM_ST.scala 32:46]
  assign _GEN_184 = 7'h3b == RADDR ? 7'h3b : _GEN_183; // @[RAM_ST.scala 32:46]
  assign _GEN_185 = 7'h3c == RADDR ? 7'h3c : _GEN_184; // @[RAM_ST.scala 32:46]
  assign _GEN_186 = 7'h3d == RADDR ? 7'h3d : _GEN_185; // @[RAM_ST.scala 32:46]
  assign _GEN_187 = 7'h3e == RADDR ? 7'h3e : _GEN_186; // @[RAM_ST.scala 32:46]
  assign _GEN_188 = 7'h3f == RADDR ? 7'h3f : _GEN_187; // @[RAM_ST.scala 32:46]
  assign _GEN_189 = 7'h40 == RADDR ? 7'h40 : _GEN_188; // @[RAM_ST.scala 32:46]
  assign _GEN_190 = 7'h41 == RADDR ? 7'h41 : _GEN_189; // @[RAM_ST.scala 32:46]
  assign _GEN_191 = 7'h42 == RADDR ? 7'h42 : _GEN_190; // @[RAM_ST.scala 32:46]
  assign _GEN_192 = 7'h43 == RADDR ? 7'h43 : _GEN_191; // @[RAM_ST.scala 32:46]
  assign _GEN_193 = 7'h44 == RADDR ? 7'h44 : _GEN_192; // @[RAM_ST.scala 32:46]
  assign _GEN_194 = 7'h45 == RADDR ? 7'h45 : _GEN_193; // @[RAM_ST.scala 32:46]
  assign _GEN_195 = 7'h46 == RADDR ? 7'h46 : _GEN_194; // @[RAM_ST.scala 32:46]
  assign _GEN_196 = 7'h47 == RADDR ? 7'h47 : _GEN_195; // @[RAM_ST.scala 32:46]
  assign _GEN_197 = 7'h48 == RADDR ? 7'h48 : _GEN_196; // @[RAM_ST.scala 32:46]
  assign _GEN_198 = 7'h49 == RADDR ? 7'h49 : _GEN_197; // @[RAM_ST.scala 32:46]
  assign _GEN_199 = 7'h4a == RADDR ? 7'h4a : _GEN_198; // @[RAM_ST.scala 32:46]
  assign _GEN_200 = 7'h4b == RADDR ? 7'h4b : _GEN_199; // @[RAM_ST.scala 32:46]
  assign _GEN_201 = 7'h4c == RADDR ? 7'h4c : _GEN_200; // @[RAM_ST.scala 32:46]
  assign _GEN_202 = 7'h4d == RADDR ? 7'h4d : _GEN_201; // @[RAM_ST.scala 32:46]
  assign _GEN_203 = 7'h4e == RADDR ? 7'h4e : _GEN_202; // @[RAM_ST.scala 32:46]
  assign _GEN_204 = 7'h4f == RADDR ? 7'h4f : _GEN_203; // @[RAM_ST.scala 32:46]
  assign _GEN_205 = 7'h50 == RADDR ? 7'h50 : _GEN_204; // @[RAM_ST.scala 32:46]
  assign _GEN_206 = 7'h51 == RADDR ? 7'h51 : _GEN_205; // @[RAM_ST.scala 32:46]
  assign _GEN_207 = 7'h52 == RADDR ? 7'h52 : _GEN_206; // @[RAM_ST.scala 32:46]
  assign _GEN_208 = 7'h53 == RADDR ? 7'h53 : _GEN_207; // @[RAM_ST.scala 32:46]
  assign _GEN_209 = 7'h54 == RADDR ? 7'h54 : _GEN_208; // @[RAM_ST.scala 32:46]
  assign _GEN_210 = 7'h55 == RADDR ? 7'h55 : _GEN_209; // @[RAM_ST.scala 32:46]
  assign _GEN_211 = 7'h56 == RADDR ? 7'h56 : _GEN_210; // @[RAM_ST.scala 32:46]
  assign _GEN_212 = 7'h57 == RADDR ? 7'h57 : _GEN_211; // @[RAM_ST.scala 32:46]
  assign _GEN_213 = 7'h58 == RADDR ? 7'h58 : _GEN_212; // @[RAM_ST.scala 32:46]
  assign _GEN_214 = 7'h59 == RADDR ? 7'h59 : _GEN_213; // @[RAM_ST.scala 32:46]
  assign _GEN_215 = 7'h5a == RADDR ? 7'h5a : _GEN_214; // @[RAM_ST.scala 32:46]
  assign _GEN_216 = 7'h5b == RADDR ? 7'h5b : _GEN_215; // @[RAM_ST.scala 32:46]
  assign _GEN_217 = 7'h5c == RADDR ? 7'h5c : _GEN_216; // @[RAM_ST.scala 32:46]
  assign _GEN_218 = 7'h5d == RADDR ? 7'h5d : _GEN_217; // @[RAM_ST.scala 32:46]
  assign _GEN_219 = 7'h5e == RADDR ? 7'h5e : _GEN_218; // @[RAM_ST.scala 32:46]
  assign _GEN_220 = 7'h5f == RADDR ? 7'h5f : _GEN_219; // @[RAM_ST.scala 32:46]
  assign _GEN_221 = 7'h60 == RADDR ? 7'h60 : _GEN_220; // @[RAM_ST.scala 32:46]
  assign _GEN_222 = 7'h61 == RADDR ? 7'h61 : _GEN_221; // @[RAM_ST.scala 32:46]
  assign _GEN_223 = 7'h62 == RADDR ? 7'h62 : _GEN_222; // @[RAM_ST.scala 32:46]
  assign _GEN_224 = 7'h63 == RADDR ? 7'h63 : _GEN_223; // @[RAM_ST.scala 32:46]
  assign _GEN_225 = 7'h64 == RADDR ? 7'h64 : _GEN_224; // @[RAM_ST.scala 32:46]
  assign _GEN_226 = 7'h65 == RADDR ? 7'h65 : _GEN_225; // @[RAM_ST.scala 32:46]
  assign _GEN_227 = 7'h66 == RADDR ? 7'h66 : _GEN_226; // @[RAM_ST.scala 32:46]
  assign _GEN_228 = 7'h67 == RADDR ? 7'h67 : _GEN_227; // @[RAM_ST.scala 32:46]
  assign _GEN_229 = 7'h68 == RADDR ? 7'h68 : _GEN_228; // @[RAM_ST.scala 32:46]
  assign _GEN_230 = 7'h69 == RADDR ? 7'h69 : _GEN_229; // @[RAM_ST.scala 32:46]
  assign _GEN_231 = 7'h6a == RADDR ? 7'h6a : _GEN_230; // @[RAM_ST.scala 32:46]
  assign _GEN_232 = 7'h6b == RADDR ? 7'h6b : _GEN_231; // @[RAM_ST.scala 32:46]
  assign _GEN_233 = 7'h6c == RADDR ? 7'h6c : _GEN_232; // @[RAM_ST.scala 32:46]
  assign _GEN_234 = 7'h6d == RADDR ? 7'h6d : _GEN_233; // @[RAM_ST.scala 32:46]
  assign _GEN_235 = 7'h6e == RADDR ? 7'h6e : _GEN_234; // @[RAM_ST.scala 32:46]
  assign _GEN_236 = 7'h6f == RADDR ? 7'h6f : _GEN_235; // @[RAM_ST.scala 32:46]
  assign _GEN_237 = 7'h70 == RADDR ? 7'h70 : _GEN_236; // @[RAM_ST.scala 32:46]
  assign _GEN_238 = 7'h71 == RADDR ? 7'h71 : _GEN_237; // @[RAM_ST.scala 32:46]
  assign _GEN_239 = 7'h72 == RADDR ? 7'h72 : _GEN_238; // @[RAM_ST.scala 32:46]
  assign _GEN_240 = 7'h73 == RADDR ? 7'h73 : _GEN_239; // @[RAM_ST.scala 32:46]
  assign _GEN_241 = 7'h74 == RADDR ? 7'h74 : _GEN_240; // @[RAM_ST.scala 32:46]
  assign _GEN_242 = 7'h75 == RADDR ? 7'h75 : _GEN_241; // @[RAM_ST.scala 32:46]
  assign _GEN_243 = 7'h76 == RADDR ? 7'h76 : _GEN_242; // @[RAM_ST.scala 32:46]
  assign _GEN_244 = 7'h77 == RADDR ? 7'h77 : _GEN_243; // @[RAM_ST.scala 32:46]
  assign _T_3 = {{1'd0}, _GEN_244}; // @[RAM_ST.scala 32:46]
  assign RDATA = ram__T_8_data; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 120; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_8_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_8_addr_pipe_0 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_2_en & ram__T_2_mask) begin
      ram[ram__T_2_addr] <= ram__T_2_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_8_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_8_addr_pipe_0 <= _T_3[6:0];
    end
  end
endmodule
module ShiftT(
  input         clock,
  input         reset,
  input         valid_up,
  input  [15:0] I,
  output [15:0] O
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_RDATA; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [15:0] RAM_ST_WDATA; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [6:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [6:0] _T_3; // @[Counter.scala 38:22]
  reg [15:0] _T_8; // @[ShiftT.scala 51:17]
  reg [31:0] _RAND_1;
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA(RAM_ST_RDATA),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA(RAM_ST_WDATA)
  );
  NestedCounters NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 7'h77; // @[Counter.scala 37:24]
  assign _T_3 = value + 7'h1; // @[Counter.scala 38:22]
  assign O = _T_8; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 7'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA = I; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_8 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 7'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 7'h0;
      end else begin
        value <= _T_3;
      end
    end
    _T_8 <= RAM_ST_RDATA;
  end
endmodule
module ShiftTS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  input  [15:0] I_8,
  input  [15:0] I_9,
  input  [15:0] I_10,
  input  [15:0] I_11,
  input  [15:0] I_12,
  input  [15:0] I_13,
  input  [15:0] I_14,
  input  [15:0] I_15,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7,
  output [15:0] O_8,
  output [15:0] O_9,
  output [15:0] O_10,
  output [15:0] O_11,
  output [15:0] O_12,
  output [15:0] O_13,
  output [15:0] O_14,
  output [15:0] O_15
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_1_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_1_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_2_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_2_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_3_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_3_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_4_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_4_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_5_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_5_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_6_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_6_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_7_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_7_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_8_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_8_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_9_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_9_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_10_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_10_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_11_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_11_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_12_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_12_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_13_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_13_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_14_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_14_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_valid_up; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_15_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_15_O; // @[ShiftTS.scala 32:34]
  reg  _T; // @[ShiftTS.scala 39:24]
  reg [31:0] _RAND_0;
  ShiftT ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I(ShiftT_I),
    .O(ShiftT_O)
  );
  ShiftT ShiftT_1 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_1_clock),
    .reset(ShiftT_1_reset),
    .valid_up(ShiftT_1_valid_up),
    .I(ShiftT_1_I),
    .O(ShiftT_1_O)
  );
  ShiftT ShiftT_2 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_2_clock),
    .reset(ShiftT_2_reset),
    .valid_up(ShiftT_2_valid_up),
    .I(ShiftT_2_I),
    .O(ShiftT_2_O)
  );
  ShiftT ShiftT_3 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_3_clock),
    .reset(ShiftT_3_reset),
    .valid_up(ShiftT_3_valid_up),
    .I(ShiftT_3_I),
    .O(ShiftT_3_O)
  );
  ShiftT ShiftT_4 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_4_clock),
    .reset(ShiftT_4_reset),
    .valid_up(ShiftT_4_valid_up),
    .I(ShiftT_4_I),
    .O(ShiftT_4_O)
  );
  ShiftT ShiftT_5 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_5_clock),
    .reset(ShiftT_5_reset),
    .valid_up(ShiftT_5_valid_up),
    .I(ShiftT_5_I),
    .O(ShiftT_5_O)
  );
  ShiftT ShiftT_6 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_6_clock),
    .reset(ShiftT_6_reset),
    .valid_up(ShiftT_6_valid_up),
    .I(ShiftT_6_I),
    .O(ShiftT_6_O)
  );
  ShiftT ShiftT_7 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_7_clock),
    .reset(ShiftT_7_reset),
    .valid_up(ShiftT_7_valid_up),
    .I(ShiftT_7_I),
    .O(ShiftT_7_O)
  );
  ShiftT ShiftT_8 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_8_clock),
    .reset(ShiftT_8_reset),
    .valid_up(ShiftT_8_valid_up),
    .I(ShiftT_8_I),
    .O(ShiftT_8_O)
  );
  ShiftT ShiftT_9 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_9_clock),
    .reset(ShiftT_9_reset),
    .valid_up(ShiftT_9_valid_up),
    .I(ShiftT_9_I),
    .O(ShiftT_9_O)
  );
  ShiftT ShiftT_10 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_10_clock),
    .reset(ShiftT_10_reset),
    .valid_up(ShiftT_10_valid_up),
    .I(ShiftT_10_I),
    .O(ShiftT_10_O)
  );
  ShiftT ShiftT_11 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_11_clock),
    .reset(ShiftT_11_reset),
    .valid_up(ShiftT_11_valid_up),
    .I(ShiftT_11_I),
    .O(ShiftT_11_O)
  );
  ShiftT ShiftT_12 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_12_clock),
    .reset(ShiftT_12_reset),
    .valid_up(ShiftT_12_valid_up),
    .I(ShiftT_12_I),
    .O(ShiftT_12_O)
  );
  ShiftT ShiftT_13 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_13_clock),
    .reset(ShiftT_13_reset),
    .valid_up(ShiftT_13_valid_up),
    .I(ShiftT_13_I),
    .O(ShiftT_13_O)
  );
  ShiftT ShiftT_14 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_14_clock),
    .reset(ShiftT_14_reset),
    .valid_up(ShiftT_14_valid_up),
    .I(ShiftT_14_I),
    .O(ShiftT_14_O)
  );
  ShiftT ShiftT_15 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_15_clock),
    .reset(ShiftT_15_reset),
    .valid_up(ShiftT_15_valid_up),
    .I(ShiftT_15_I),
    .O(ShiftT_15_O)
  );
  assign valid_down = _T; // @[ShiftTS.scala 39:14]
  assign O_0 = ShiftT_O; // @[ShiftTS.scala 34:36]
  assign O_1 = ShiftT_1_O; // @[ShiftTS.scala 34:36]
  assign O_2 = ShiftT_2_O; // @[ShiftTS.scala 34:36]
  assign O_3 = ShiftT_3_O; // @[ShiftTS.scala 34:36]
  assign O_4 = ShiftT_4_O; // @[ShiftTS.scala 34:36]
  assign O_5 = ShiftT_5_O; // @[ShiftTS.scala 34:36]
  assign O_6 = ShiftT_6_O; // @[ShiftTS.scala 34:36]
  assign O_7 = ShiftT_7_O; // @[ShiftTS.scala 34:36]
  assign O_8 = ShiftT_8_O; // @[ShiftTS.scala 34:36]
  assign O_9 = ShiftT_9_O; // @[ShiftTS.scala 34:36]
  assign O_10 = ShiftT_10_O; // @[ShiftTS.scala 34:36]
  assign O_11 = ShiftT_11_O; // @[ShiftTS.scala 34:36]
  assign O_12 = ShiftT_12_O; // @[ShiftTS.scala 34:36]
  assign O_13 = ShiftT_13_O; // @[ShiftTS.scala 34:36]
  assign O_14 = ShiftT_14_O; // @[ShiftTS.scala 34:36]
  assign O_15 = ShiftT_15_O; // @[ShiftTS.scala 34:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_I = I_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_1_clock = clock;
  assign ShiftT_1_reset = reset;
  assign ShiftT_1_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_1_I = I_1; // @[ShiftTS.scala 33:24]
  assign ShiftT_2_clock = clock;
  assign ShiftT_2_reset = reset;
  assign ShiftT_2_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_2_I = I_2; // @[ShiftTS.scala 33:24]
  assign ShiftT_3_clock = clock;
  assign ShiftT_3_reset = reset;
  assign ShiftT_3_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_3_I = I_3; // @[ShiftTS.scala 33:24]
  assign ShiftT_4_clock = clock;
  assign ShiftT_4_reset = reset;
  assign ShiftT_4_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_4_I = I_4; // @[ShiftTS.scala 33:24]
  assign ShiftT_5_clock = clock;
  assign ShiftT_5_reset = reset;
  assign ShiftT_5_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_5_I = I_5; // @[ShiftTS.scala 33:24]
  assign ShiftT_6_clock = clock;
  assign ShiftT_6_reset = reset;
  assign ShiftT_6_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_6_I = I_6; // @[ShiftTS.scala 33:24]
  assign ShiftT_7_clock = clock;
  assign ShiftT_7_reset = reset;
  assign ShiftT_7_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_7_I = I_7; // @[ShiftTS.scala 33:24]
  assign ShiftT_8_clock = clock;
  assign ShiftT_8_reset = reset;
  assign ShiftT_8_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_8_I = I_8; // @[ShiftTS.scala 33:24]
  assign ShiftT_9_clock = clock;
  assign ShiftT_9_reset = reset;
  assign ShiftT_9_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_9_I = I_9; // @[ShiftTS.scala 33:24]
  assign ShiftT_10_clock = clock;
  assign ShiftT_10_reset = reset;
  assign ShiftT_10_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_10_I = I_10; // @[ShiftTS.scala 33:24]
  assign ShiftT_11_clock = clock;
  assign ShiftT_11_reset = reset;
  assign ShiftT_11_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_11_I = I_11; // @[ShiftTS.scala 33:24]
  assign ShiftT_12_clock = clock;
  assign ShiftT_12_reset = reset;
  assign ShiftT_12_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_12_I = I_12; // @[ShiftTS.scala 33:24]
  assign ShiftT_13_clock = clock;
  assign ShiftT_13_reset = reset;
  assign ShiftT_13_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_13_I = I_13; // @[ShiftTS.scala 33:24]
  assign ShiftT_14_clock = clock;
  assign ShiftT_14_reset = reset;
  assign ShiftT_14_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_14_I = I_14; // @[ShiftTS.scala 33:24]
  assign ShiftT_15_clock = clock;
  assign ShiftT_15_reset = reset;
  assign ShiftT_15_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_15_I = I_15; // @[ShiftTS.scala 33:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 1'h0;
    end else begin
      _T <= valid_up;
    end
  end
endmodule
module ShiftT_32(
  input         clock,
  input  [15:0] I,
  output [15:0] O
);
  reg [15:0] _T; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O = _T; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= I;
  end
endmodule
module ShiftTS_2(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  input  [15:0] I_8,
  input  [15:0] I_9,
  input  [15:0] I_10,
  input  [15:0] I_11,
  input  [15:0] I_12,
  input  [15:0] I_13,
  input  [15:0] I_14,
  input  [15:0] I_15,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7,
  output [15:0] O_8,
  output [15:0] O_9,
  output [15:0] O_10,
  output [15:0] O_11,
  output [15:0] O_12,
  output [15:0] O_13,
  output [15:0] O_14,
  output [15:0] O_15
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_I; // @[ShiftTS.scala 32:34]
  wire [15:0] ShiftT_O; // @[ShiftTS.scala 32:34]
  reg  _T; // @[ShiftTS.scala 39:24]
  reg [31:0] _RAND_0;
  ShiftT_32 ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .I(ShiftT_I),
    .O(ShiftT_O)
  );
  assign valid_down = _T; // @[ShiftTS.scala 39:14]
  assign O_0 = ShiftT_O; // @[ShiftTS.scala 34:36]
  assign O_1 = I_0; // @[ShiftTS.scala 29:36]
  assign O_2 = I_1; // @[ShiftTS.scala 29:36]
  assign O_3 = I_2; // @[ShiftTS.scala 29:36]
  assign O_4 = I_3; // @[ShiftTS.scala 29:36]
  assign O_5 = I_4; // @[ShiftTS.scala 29:36]
  assign O_6 = I_5; // @[ShiftTS.scala 29:36]
  assign O_7 = I_6; // @[ShiftTS.scala 29:36]
  assign O_8 = I_7; // @[ShiftTS.scala 29:36]
  assign O_9 = I_8; // @[ShiftTS.scala 29:36]
  assign O_10 = I_9; // @[ShiftTS.scala 29:36]
  assign O_11 = I_10; // @[ShiftTS.scala 29:36]
  assign O_12 = I_11; // @[ShiftTS.scala 29:36]
  assign O_13 = I_12; // @[ShiftTS.scala 29:36]
  assign O_14 = I_13; // @[ShiftTS.scala 29:36]
  assign O_15 = I_14; // @[ShiftTS.scala 29:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I = I_15; // @[ShiftTS.scala 33:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 1'h0;
    end else begin
      _T <= valid_up;
    end
  end
endmodule
module SSeqTupleCreator(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  input  [15:0] I1,
  output [15:0] O_0,
  output [15:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I0_3,
  input  [15:0] I0_4,
  input  [15:0] I0_5,
  input  [15:0] I0_6,
  input  [15:0] I0_7,
  input  [15:0] I0_8,
  input  [15:0] I0_9,
  input  [15:0] I0_10,
  input  [15:0] I0_11,
  input  [15:0] I0_12,
  input  [15:0] I0_13,
  input  [15:0] I0_14,
  input  [15:0] I0_15,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  input  [15:0] I1_8,
  input  [15:0] I1_9,
  input  [15:0] I1_10,
  input  [15:0] I1_11,
  input  [15:0] I1_12,
  input  [15:0] I1_13,
  input  [15:0] I1_14,
  input  [15:0] I1_15,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_15_0,
  output [15:0] O_15_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  SSeqTupleCreator other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  SSeqTupleCreator other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  SSeqTupleCreator other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1)
  );
  SSeqTupleCreator other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1)
  );
  SSeqTupleCreator other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1)
  );
  SSeqTupleCreator other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1)
  );
  SSeqTupleCreator other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0(other_ops_7_I0),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1)
  );
  SSeqTupleCreator other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0(other_ops_8_I0),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1)
  );
  SSeqTupleCreator other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0(other_ops_9_I0),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1)
  );
  SSeqTupleCreator other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0(other_ops_10_I0),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1)
  );
  SSeqTupleCreator other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0(other_ops_11_I0),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1)
  );
  SSeqTupleCreator other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0(other_ops_12_I0),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1)
  );
  SSeqTupleCreator other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0(other_ops_13_I0),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1)
  );
  SSeqTupleCreator other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0(other_ops_14_I0),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0 = I0_8; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0 = I0_9; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0 = I0_10; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0 = I0_11; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0 = I0_12; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0 = I0_13; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0 = I0_14; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0 = I0_15; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I0_3,
  input  [15:0] I0_4,
  input  [15:0] I0_5,
  input  [15:0] I0_6,
  input  [15:0] I0_7,
  input  [15:0] I0_8,
  input  [15:0] I0_9,
  input  [15:0] I0_10,
  input  [15:0] I0_11,
  input  [15:0] I0_12,
  input  [15:0] I0_13,
  input  [15:0] I0_14,
  input  [15:0] I0_15,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  input  [15:0] I1_8,
  input  [15:0] I1_9,
  input  [15:0] I1_10,
  input  [15:0] I1_11,
  input  [15:0] I1_12,
  input  [15:0] I1_13,
  input  [15:0] I1_14,
  input  [15:0] I1_15,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_15_0,
  output [15:0] O_15_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I0_8(op_I0_8),
    .I0_9(op_I0_9),
    .I0_10(op_I0_10),
    .I0_11(op_I0_11),
    .I0_12(op_I0_12),
    .I0_13(op_I0_13),
    .I0_14(op_I0_14),
    .I0_15(op_I0_15),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .I1_8(op_I1_8),
    .I1_9(op_I1_9),
    .I1_10(op_I1_10),
    .I1_11(op_I1_11),
    .I1_12(op_I1_12),
    .I1_13(op_I1_13),
    .I1_14(op_I1_14),
    .I1_15(op_I1_15),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_8_0 = op_O_8_0; // @[Map2T.scala 17:7]
  assign O_8_1 = op_O_8_1; // @[Map2T.scala 17:7]
  assign O_9_0 = op_O_9_0; // @[Map2T.scala 17:7]
  assign O_9_1 = op_O_9_1; // @[Map2T.scala 17:7]
  assign O_10_0 = op_O_10_0; // @[Map2T.scala 17:7]
  assign O_10_1 = op_O_10_1; // @[Map2T.scala 17:7]
  assign O_11_0 = op_O_11_0; // @[Map2T.scala 17:7]
  assign O_11_1 = op_O_11_1; // @[Map2T.scala 17:7]
  assign O_12_0 = op_O_12_0; // @[Map2T.scala 17:7]
  assign O_12_1 = op_O_12_1; // @[Map2T.scala 17:7]
  assign O_13_0 = op_O_13_0; // @[Map2T.scala 17:7]
  assign O_13_1 = op_O_13_1; // @[Map2T.scala 17:7]
  assign O_14_0 = op_O_14_0; // @[Map2T.scala 17:7]
  assign O_14_1 = op_O_14_1; // @[Map2T.scala 17:7]
  assign O_15_0 = op_O_15_0; // @[Map2T.scala 17:7]
  assign O_15_1 = op_O_15_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I0_8 = I0_8; // @[Map2T.scala 15:11]
  assign op_I0_9 = I0_9; // @[Map2T.scala 15:11]
  assign op_I0_10 = I0_10; // @[Map2T.scala 15:11]
  assign op_I0_11 = I0_11; // @[Map2T.scala 15:11]
  assign op_I0_12 = I0_12; // @[Map2T.scala 15:11]
  assign op_I0_13 = I0_13; // @[Map2T.scala 15:11]
  assign op_I0_14 = I0_14; // @[Map2T.scala 15:11]
  assign op_I0_15 = I0_15; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
  assign op_I1_8 = I1_8; // @[Map2T.scala 16:11]
  assign op_I1_9 = I1_9; // @[Map2T.scala 16:11]
  assign op_I1_10 = I1_10; // @[Map2T.scala 16:11]
  assign op_I1_11 = I1_11; // @[Map2T.scala 16:11]
  assign op_I1_12 = I1_12; // @[Map2T.scala 16:11]
  assign op_I1_13 = I1_13; // @[Map2T.scala 16:11]
  assign op_I1_14 = I1_14; // @[Map2T.scala 16:11]
  assign op_I1_15 = I1_15; // @[Map2T.scala 16:11]
endmodule
module FIFO_2(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  input  [15:0] I_8,
  input  [15:0] I_9,
  input  [15:0] I_10,
  input  [15:0] I_11,
  input  [15:0] I_12,
  input  [15:0] I_13,
  input  [15:0] I_14,
  input  [15:0] I_15,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7,
  output [15:0] O_8,
  output [15:0] O_9,
  output [15:0] O_10,
  output [15:0] O_11,
  output [15:0] O_12,
  output [15:0] O_13,
  output [15:0] O_14,
  output [15:0] O_15
);
  reg [15:0] _T__0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [15:0] _T__0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [15:0] _T__0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__0__T_17_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T__0__T_17_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [15:0] _T__1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_4;
  wire [15:0] _T__1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_5;
  wire [15:0] _T__1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__1__T_17_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [1:0] _T__1__T_17_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [15:0] _T__2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_8;
  wire [15:0] _T__2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_9;
  wire [15:0] _T__2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__2__T_17_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [1:0] _T__2__T_17_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [15:0] _T__3 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_12;
  wire [15:0] _T__3__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_13;
  wire [15:0] _T__3__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__3__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__3__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__3__T_17_en_pipe_0;
  reg [31:0] _RAND_14;
  reg [1:0] _T__3__T_17_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [15:0] _T__4 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_16;
  wire [15:0] _T__4__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_17;
  wire [15:0] _T__4__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__4__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__4__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__4__T_17_en_pipe_0;
  reg [31:0] _RAND_18;
  reg [1:0] _T__4__T_17_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [15:0] _T__5 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_20;
  wire [15:0] _T__5__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_21;
  wire [15:0] _T__5__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__5__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__5__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__5__T_17_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [1:0] _T__5__T_17_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [15:0] _T__6 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_24;
  wire [15:0] _T__6__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_25;
  wire [15:0] _T__6__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__6__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__6__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__6__T_17_en_pipe_0;
  reg [31:0] _RAND_26;
  reg [1:0] _T__6__T_17_addr_pipe_0;
  reg [31:0] _RAND_27;
  reg [15:0] _T__7 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_28;
  wire [15:0] _T__7__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_29;
  wire [15:0] _T__7__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__7__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__7__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__7__T_17_en_pipe_0;
  reg [31:0] _RAND_30;
  reg [1:0] _T__7__T_17_addr_pipe_0;
  reg [31:0] _RAND_31;
  reg [15:0] _T__8 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_32;
  wire [15:0] _T__8__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_33;
  wire [15:0] _T__8__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__8__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__8__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__8__T_17_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [1:0] _T__8__T_17_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [15:0] _T__9 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_36;
  wire [15:0] _T__9__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_37;
  wire [15:0] _T__9__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__9__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__9__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__9__T_17_en_pipe_0;
  reg [31:0] _RAND_38;
  reg [1:0] _T__9__T_17_addr_pipe_0;
  reg [31:0] _RAND_39;
  reg [15:0] _T__10 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_40;
  wire [15:0] _T__10__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_41;
  wire [15:0] _T__10__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__10__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__10__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__10__T_17_en_pipe_0;
  reg [31:0] _RAND_42;
  reg [1:0] _T__10__T_17_addr_pipe_0;
  reg [31:0] _RAND_43;
  reg [15:0] _T__11 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_44;
  wire [15:0] _T__11__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_45;
  wire [15:0] _T__11__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__11__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__11__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__11__T_17_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [1:0] _T__11__T_17_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [15:0] _T__12 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_48;
  wire [15:0] _T__12__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_49;
  wire [15:0] _T__12__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__12__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__12__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__12__T_17_en_pipe_0;
  reg [31:0] _RAND_50;
  reg [1:0] _T__12__T_17_addr_pipe_0;
  reg [31:0] _RAND_51;
  reg [15:0] _T__13 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_52;
  wire [15:0] _T__13__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_53;
  wire [15:0] _T__13__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__13__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__13__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__13__T_17_en_pipe_0;
  reg [31:0] _RAND_54;
  reg [1:0] _T__13__T_17_addr_pipe_0;
  reg [31:0] _RAND_55;
  reg [15:0] _T__14 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_56;
  wire [15:0] _T__14__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_57;
  wire [15:0] _T__14__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__14__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__14__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__14__T_17_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [1:0] _T__14__T_17_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [15:0] _T__15 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_60;
  wire [15:0] _T__15__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_61;
  wire [15:0] _T__15__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__15__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__15__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__15__T_17_en_pipe_0;
  reg [31:0] _RAND_62;
  reg [1:0] _T__15__T_17_addr_pipe_0;
  reg [31:0] _RAND_63;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_64;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_65;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_66;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_11; // @[Counter.scala 38:22]
  wire  _T_12; // @[FIFO.scala 42:39]
  wire  _T_18; // @[Counter.scala 37:24]
  wire [1:0] _T_20; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  wire  _GEN_70; // @[FIFO.scala 39:15]
  assign _T__0__T_17_addr = _T__0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0__T_17_data = _T__0[_T__0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__0__T_17_data = _T__0__T_17_addr >= 2'h3 ? _RAND_1[15:0] : _T__0[_T__0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0__T_5_data = I_0;
  assign _T__0__T_5_addr = value_2;
  assign _T__0__T_5_mask = 1'h1;
  assign _T__0__T_5_en = valid_up;
  assign _T__1__T_17_addr = _T__1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1__T_17_data = _T__1[_T__1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__1__T_17_data = _T__1__T_17_addr >= 2'h3 ? _RAND_5[15:0] : _T__1[_T__1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1__T_5_data = I_1;
  assign _T__1__T_5_addr = value_2;
  assign _T__1__T_5_mask = 1'h1;
  assign _T__1__T_5_en = valid_up;
  assign _T__2__T_17_addr = _T__2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2__T_17_data = _T__2[_T__2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__2__T_17_data = _T__2__T_17_addr >= 2'h3 ? _RAND_9[15:0] : _T__2[_T__2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2__T_5_data = I_2;
  assign _T__2__T_5_addr = value_2;
  assign _T__2__T_5_mask = 1'h1;
  assign _T__2__T_5_en = valid_up;
  assign _T__3__T_17_addr = _T__3__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3__T_17_data = _T__3[_T__3__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__3__T_17_data = _T__3__T_17_addr >= 2'h3 ? _RAND_13[15:0] : _T__3[_T__3__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3__T_5_data = I_3;
  assign _T__3__T_5_addr = value_2;
  assign _T__3__T_5_mask = 1'h1;
  assign _T__3__T_5_en = valid_up;
  assign _T__4__T_17_addr = _T__4__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4__T_17_data = _T__4[_T__4__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__4__T_17_data = _T__4__T_17_addr >= 2'h3 ? _RAND_17[15:0] : _T__4[_T__4__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4__T_5_data = I_4;
  assign _T__4__T_5_addr = value_2;
  assign _T__4__T_5_mask = 1'h1;
  assign _T__4__T_5_en = valid_up;
  assign _T__5__T_17_addr = _T__5__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5__T_17_data = _T__5[_T__5__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__5__T_17_data = _T__5__T_17_addr >= 2'h3 ? _RAND_21[15:0] : _T__5[_T__5__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5__T_5_data = I_5;
  assign _T__5__T_5_addr = value_2;
  assign _T__5__T_5_mask = 1'h1;
  assign _T__5__T_5_en = valid_up;
  assign _T__6__T_17_addr = _T__6__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6__T_17_data = _T__6[_T__6__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__6__T_17_data = _T__6__T_17_addr >= 2'h3 ? _RAND_25[15:0] : _T__6[_T__6__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6__T_5_data = I_6;
  assign _T__6__T_5_addr = value_2;
  assign _T__6__T_5_mask = 1'h1;
  assign _T__6__T_5_en = valid_up;
  assign _T__7__T_17_addr = _T__7__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7__T_17_data = _T__7[_T__7__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__7__T_17_data = _T__7__T_17_addr >= 2'h3 ? _RAND_29[15:0] : _T__7[_T__7__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7__T_5_data = I_7;
  assign _T__7__T_5_addr = value_2;
  assign _T__7__T_5_mask = 1'h1;
  assign _T__7__T_5_en = valid_up;
  assign _T__8__T_17_addr = _T__8__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8__T_17_data = _T__8[_T__8__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__8__T_17_data = _T__8__T_17_addr >= 2'h3 ? _RAND_33[15:0] : _T__8[_T__8__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8__T_5_data = I_8;
  assign _T__8__T_5_addr = value_2;
  assign _T__8__T_5_mask = 1'h1;
  assign _T__8__T_5_en = valid_up;
  assign _T__9__T_17_addr = _T__9__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9__T_17_data = _T__9[_T__9__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__9__T_17_data = _T__9__T_17_addr >= 2'h3 ? _RAND_37[15:0] : _T__9[_T__9__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9__T_5_data = I_9;
  assign _T__9__T_5_addr = value_2;
  assign _T__9__T_5_mask = 1'h1;
  assign _T__9__T_5_en = valid_up;
  assign _T__10__T_17_addr = _T__10__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10__T_17_data = _T__10[_T__10__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__10__T_17_data = _T__10__T_17_addr >= 2'h3 ? _RAND_41[15:0] : _T__10[_T__10__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10__T_5_data = I_10;
  assign _T__10__T_5_addr = value_2;
  assign _T__10__T_5_mask = 1'h1;
  assign _T__10__T_5_en = valid_up;
  assign _T__11__T_17_addr = _T__11__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11__T_17_data = _T__11[_T__11__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__11__T_17_data = _T__11__T_17_addr >= 2'h3 ? _RAND_45[15:0] : _T__11[_T__11__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11__T_5_data = I_11;
  assign _T__11__T_5_addr = value_2;
  assign _T__11__T_5_mask = 1'h1;
  assign _T__11__T_5_en = valid_up;
  assign _T__12__T_17_addr = _T__12__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12__T_17_data = _T__12[_T__12__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__12__T_17_data = _T__12__T_17_addr >= 2'h3 ? _RAND_49[15:0] : _T__12[_T__12__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12__T_5_data = I_12;
  assign _T__12__T_5_addr = value_2;
  assign _T__12__T_5_mask = 1'h1;
  assign _T__12__T_5_en = valid_up;
  assign _T__13__T_17_addr = _T__13__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13__T_17_data = _T__13[_T__13__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__13__T_17_data = _T__13__T_17_addr >= 2'h3 ? _RAND_53[15:0] : _T__13[_T__13__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13__T_5_data = I_13;
  assign _T__13__T_5_addr = value_2;
  assign _T__13__T_5_mask = 1'h1;
  assign _T__13__T_5_en = valid_up;
  assign _T__14__T_17_addr = _T__14__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14__T_17_data = _T__14[_T__14__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__14__T_17_data = _T__14__T_17_addr >= 2'h3 ? _RAND_57[15:0] : _T__14[_T__14__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14__T_5_data = I_14;
  assign _T__14__T_5_addr = value_2;
  assign _T__14__T_5_mask = 1'h1;
  assign _T__14__T_5_en = valid_up;
  assign _T__15__T_17_addr = _T__15__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15__T_17_data = _T__15[_T__15__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__15__T_17_data = _T__15__T_17_addr >= 2'h3 ? _RAND_61[15:0] : _T__15[_T__15__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15__T_5_data = I_15;
  assign _T__15__T_5_addr = value_2;
  assign _T__15__T_5_mask = 1'h1;
  assign _T__15__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_11 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_12 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_18 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_20 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_12 & _T_12; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0 = _T__0__T_17_data; // @[FIFO.scala 43:11]
  assign O_1 = _T__1__T_17_data; // @[FIFO.scala 43:11]
  assign O_2 = _T__2__T_17_data; // @[FIFO.scala 43:11]
  assign O_3 = _T__3__T_17_data; // @[FIFO.scala 43:11]
  assign O_4 = _T__4__T_17_data; // @[FIFO.scala 43:11]
  assign O_5 = _T__5__T_17_data; // @[FIFO.scala 43:11]
  assign O_6 = _T__6__T_17_data; // @[FIFO.scala 43:11]
  assign O_7 = _T__7__T_17_data; // @[FIFO.scala 43:11]
  assign O_8 = _T__8__T_17_data; // @[FIFO.scala 43:11]
  assign O_9 = _T__9__T_17_data; // @[FIFO.scala 43:11]
  assign O_10 = _T__10__T_17_data; // @[FIFO.scala 43:11]
  assign O_11 = _T__11__T_17_data; // @[FIFO.scala 43:11]
  assign O_12 = _T__12__T_17_data; // @[FIFO.scala 43:11]
  assign O_13 = _T__13__T_17_data; // @[FIFO.scala 43:11]
  assign O_14 = _T__14__T_17_data; // @[FIFO.scala 43:11]
  assign O_15 = _T__15__T_17_data; // @[FIFO.scala 43:11]
  assign _GEN_70 = valid_up & _T_6; // @[FIFO.scala 39:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__0[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0__T_17_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__0__T_17_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__1[initvar] = _RAND_4[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__1__T_17_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__1__T_17_addr_pipe_0 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__2[initvar] = _RAND_8[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__2__T_17_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__2__T_17_addr_pipe_0 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__3[initvar] = _RAND_12[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__3__T_17_en_pipe_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__3__T_17_addr_pipe_0 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__4[initvar] = _RAND_16[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__4__T_17_en_pipe_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__4__T_17_addr_pipe_0 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__5[initvar] = _RAND_20[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__5__T_17_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__5__T_17_addr_pipe_0 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__6[initvar] = _RAND_24[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__6__T_17_en_pipe_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__6__T_17_addr_pipe_0 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__7[initvar] = _RAND_28[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__7__T_17_en_pipe_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__7__T_17_addr_pipe_0 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__8[initvar] = _RAND_32[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__8__T_17_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__8__T_17_addr_pipe_0 = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__9[initvar] = _RAND_36[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_37 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__9__T_17_en_pipe_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__9__T_17_addr_pipe_0 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__10[initvar] = _RAND_40[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_41 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T__10__T_17_en_pipe_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T__10__T_17_addr_pipe_0 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__11[initvar] = _RAND_44[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T__11__T_17_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T__11__T_17_addr_pipe_0 = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__12[initvar] = _RAND_48[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_49 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T__12__T_17_en_pipe_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T__12__T_17_addr_pipe_0 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__13[initvar] = _RAND_52[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_53 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T__13__T_17_en_pipe_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T__13__T_17_addr_pipe_0 = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__14[initvar] = _RAND_56[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T__14__T_17_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T__14__T_17_addr_pipe_0 = _RAND_59[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__15[initvar] = _RAND_60[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_61 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T__15__T_17_en_pipe_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T__15__T_17_addr_pipe_0 = _RAND_63[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  value = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  value_1 = _RAND_65[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  value_2 = _RAND_66[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__0__T_5_en & _T__0__T_5_mask) begin
      _T__0[_T__0__T_5_addr] <= _T__0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__1__T_5_en & _T__1__T_5_mask) begin
      _T__1[_T__1__T_5_addr] <= _T__1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__2__T_5_en & _T__2__T_5_mask) begin
      _T__2[_T__2__T_5_addr] <= _T__2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__3__T_5_en & _T__3__T_5_mask) begin
      _T__3[_T__3__T_5_addr] <= _T__3__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__3__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__3__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__4__T_5_en & _T__4__T_5_mask) begin
      _T__4[_T__4__T_5_addr] <= _T__4__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__4__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__4__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__5__T_5_en & _T__5__T_5_mask) begin
      _T__5[_T__5__T_5_addr] <= _T__5__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__5__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__5__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__6__T_5_en & _T__6__T_5_mask) begin
      _T__6[_T__6__T_5_addr] <= _T__6__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__6__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__6__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__7__T_5_en & _T__7__T_5_mask) begin
      _T__7[_T__7__T_5_addr] <= _T__7__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__7__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__7__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__8__T_5_en & _T__8__T_5_mask) begin
      _T__8[_T__8__T_5_addr] <= _T__8__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__8__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__8__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__9__T_5_en & _T__9__T_5_mask) begin
      _T__9[_T__9__T_5_addr] <= _T__9__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__9__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__9__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__10__T_5_en & _T__10__T_5_mask) begin
      _T__10[_T__10__T_5_addr] <= _T__10__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__10__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__10__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__11__T_5_en & _T__11__T_5_mask) begin
      _T__11[_T__11__T_5_addr] <= _T__11__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__11__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__11__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__12__T_5_en & _T__12__T_5_mask) begin
      _T__12[_T__12__T_5_addr] <= _T__12__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__12__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__12__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__13__T_5_en & _T__13__T_5_mask) begin
      _T__13[_T__13__T_5_addr] <= _T__13__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__13__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__13__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__14__T_5_en & _T__14__T_5_mask) begin
      _T__14[_T__14__T_5_addr] <= _T__14__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__14__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__14__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__15__T_5_en & _T__15__T_5_mask) begin
      _T__15[_T__15__T_5_addr] <= _T__15__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__15__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__15__T_17_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_11;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_12) begin
        if (_T_18) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_20;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_70 & ~reset) begin
          $fwrite(32'h80000002,"idc inc\n"); // @[FIFO.scala 39:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SSeqTupleAppender(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I1,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I0_8_0,
  input  [15:0] I0_8_1,
  input  [15:0] I0_9_0,
  input  [15:0] I0_9_1,
  input  [15:0] I0_10_0,
  input  [15:0] I0_10_1,
  input  [15:0] I0_11_0,
  input  [15:0] I0_11_1,
  input  [15:0] I0_12_0,
  input  [15:0] I0_12_1,
  input  [15:0] I0_13_0,
  input  [15:0] I0_13_1,
  input  [15:0] I0_14_0,
  input  [15:0] I0_14_1,
  input  [15:0] I0_15_0,
  input  [15:0] I0_15_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  input  [15:0] I1_8,
  input  [15:0] I1_9,
  input  [15:0] I1_10,
  input  [15:0] I1_11,
  input  [15:0] I1_12,
  input  [15:0] I1_13,
  input  [15:0] I1_14,
  input  [15:0] I1_15,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_8_2,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_9_2,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_10_2,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_11_2,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_12_2,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_13_2,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_14_2,
  output [15:0] O_15_0,
  output [15:0] O_15_1,
  output [15:0] O_15_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  SSeqTupleAppender other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  SSeqTupleAppender other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  SSeqTupleAppender other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  SSeqTupleAppender other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  SSeqTupleAppender other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  SSeqTupleAppender other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  SSeqTupleAppender other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  SSeqTupleAppender other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  SSeqTupleAppender other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  SSeqTupleAppender other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  SSeqTupleAppender other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  SSeqTupleAppender other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  SSeqTupleAppender other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  SSeqTupleAppender other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_2_2 = other_ops_1_O_2; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_3_2 = other_ops_2_O_2; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_4_2 = other_ops_3_O_2; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_5_2 = other_ops_4_O_2; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_6_2 = other_ops_5_O_2; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_7_2 = other_ops_6_O_2; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_8_2 = other_ops_7_O_2; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_9_2 = other_ops_8_O_2; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_10_2 = other_ops_9_O_2; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_11_2 = other_ops_10_O_2; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_12_2 = other_ops_11_O_2; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_13_2 = other_ops_12_O_2; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_14_2 = other_ops_13_O_2; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign O_15_2 = other_ops_14_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I0_8_0,
  input  [15:0] I0_8_1,
  input  [15:0] I0_9_0,
  input  [15:0] I0_9_1,
  input  [15:0] I0_10_0,
  input  [15:0] I0_10_1,
  input  [15:0] I0_11_0,
  input  [15:0] I0_11_1,
  input  [15:0] I0_12_0,
  input  [15:0] I0_12_1,
  input  [15:0] I0_13_0,
  input  [15:0] I0_13_1,
  input  [15:0] I0_14_0,
  input  [15:0] I0_14_1,
  input  [15:0] I0_15_0,
  input  [15:0] I0_15_1,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  input  [15:0] I1_3,
  input  [15:0] I1_4,
  input  [15:0] I1_5,
  input  [15:0] I1_6,
  input  [15:0] I1_7,
  input  [15:0] I1_8,
  input  [15:0] I1_9,
  input  [15:0] I1_10,
  input  [15:0] I1_11,
  input  [15:0] I1_12,
  input  [15:0] I1_13,
  input  [15:0] I1_14,
  input  [15:0] I1_15,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_8_2,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_9_2,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_10_2,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_11_2,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_12_2,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_13_2,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_14_2,
  output [15:0] O_15_0,
  output [15:0] O_15_1,
  output [15:0] O_15_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_8_0(op_I0_8_0),
    .I0_8_1(op_I0_8_1),
    .I0_9_0(op_I0_9_0),
    .I0_9_1(op_I0_9_1),
    .I0_10_0(op_I0_10_0),
    .I0_10_1(op_I0_10_1),
    .I0_11_0(op_I0_11_0),
    .I0_11_1(op_I0_11_1),
    .I0_12_0(op_I0_12_0),
    .I0_12_1(op_I0_12_1),
    .I0_13_0(op_I0_13_0),
    .I0_13_1(op_I0_13_1),
    .I0_14_0(op_I0_14_0),
    .I0_14_1(op_I0_14_1),
    .I0_15_0(op_I0_15_0),
    .I0_15_1(op_I0_15_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .I1_8(op_I1_8),
    .I1_9(op_I1_9),
    .I1_10(op_I1_10),
    .I1_11(op_I1_11),
    .I1_12(op_I1_12),
    .I1_13(op_I1_13),
    .I1_14(op_I1_14),
    .I1_15(op_I1_15),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_8_2(op_O_8_2),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_9_2(op_O_9_2),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_10_2(op_O_10_2),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_11_2(op_O_11_2),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_12_2(op_O_12_2),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_13_2(op_O_13_2),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_14_2(op_O_14_2),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1),
    .O_15_2(op_O_15_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_1_2 = op_O_1_2; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_2_2 = op_O_2_2; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_3_2 = op_O_3_2; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_4_2 = op_O_4_2; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_5_2 = op_O_5_2; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_6_2 = op_O_6_2; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_7_2 = op_O_7_2; // @[Map2T.scala 17:7]
  assign O_8_0 = op_O_8_0; // @[Map2T.scala 17:7]
  assign O_8_1 = op_O_8_1; // @[Map2T.scala 17:7]
  assign O_8_2 = op_O_8_2; // @[Map2T.scala 17:7]
  assign O_9_0 = op_O_9_0; // @[Map2T.scala 17:7]
  assign O_9_1 = op_O_9_1; // @[Map2T.scala 17:7]
  assign O_9_2 = op_O_9_2; // @[Map2T.scala 17:7]
  assign O_10_0 = op_O_10_0; // @[Map2T.scala 17:7]
  assign O_10_1 = op_O_10_1; // @[Map2T.scala 17:7]
  assign O_10_2 = op_O_10_2; // @[Map2T.scala 17:7]
  assign O_11_0 = op_O_11_0; // @[Map2T.scala 17:7]
  assign O_11_1 = op_O_11_1; // @[Map2T.scala 17:7]
  assign O_11_2 = op_O_11_2; // @[Map2T.scala 17:7]
  assign O_12_0 = op_O_12_0; // @[Map2T.scala 17:7]
  assign O_12_1 = op_O_12_1; // @[Map2T.scala 17:7]
  assign O_12_2 = op_O_12_2; // @[Map2T.scala 17:7]
  assign O_13_0 = op_O_13_0; // @[Map2T.scala 17:7]
  assign O_13_1 = op_O_13_1; // @[Map2T.scala 17:7]
  assign O_13_2 = op_O_13_2; // @[Map2T.scala 17:7]
  assign O_14_0 = op_O_14_0; // @[Map2T.scala 17:7]
  assign O_14_1 = op_O_14_1; // @[Map2T.scala 17:7]
  assign O_14_2 = op_O_14_2; // @[Map2T.scala 17:7]
  assign O_15_0 = op_O_15_0; // @[Map2T.scala 17:7]
  assign O_15_1 = op_O_15_1; // @[Map2T.scala 17:7]
  assign O_15_2 = op_O_15_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0 = I0_8_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1 = I0_8_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0 = I0_9_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1 = I0_9_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0 = I0_10_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1 = I0_10_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0 = I0_11_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1 = I0_11_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0 = I0_12_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1 = I0_12_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0 = I0_13_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1 = I0_13_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0 = I0_14_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1 = I0_14_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0 = I0_15_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1 = I0_15_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
  assign op_I1_8 = I1_8; // @[Map2T.scala 16:11]
  assign op_I1_9 = I1_9; // @[Map2T.scala 16:11]
  assign op_I1_10 = I1_10; // @[Map2T.scala 16:11]
  assign op_I1_11 = I1_11; // @[Map2T.scala 16:11]
  assign op_I1_12 = I1_12; // @[Map2T.scala 16:11]
  assign op_I1_13 = I1_13; // @[Map2T.scala 16:11]
  assign op_I1_14 = I1_14; // @[Map2T.scala 16:11]
  assign op_I1_15 = I1_15; // @[Map2T.scala 16:11]
endmodule
module PartitionS(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  input  [15:0] I_4_0,
  input  [15:0] I_4_1,
  input  [15:0] I_4_2,
  input  [15:0] I_5_0,
  input  [15:0] I_5_1,
  input  [15:0] I_5_2,
  input  [15:0] I_6_0,
  input  [15:0] I_6_1,
  input  [15:0] I_6_2,
  input  [15:0] I_7_0,
  input  [15:0] I_7_1,
  input  [15:0] I_7_2,
  input  [15:0] I_8_0,
  input  [15:0] I_8_1,
  input  [15:0] I_8_2,
  input  [15:0] I_9_0,
  input  [15:0] I_9_1,
  input  [15:0] I_9_2,
  input  [15:0] I_10_0,
  input  [15:0] I_10_1,
  input  [15:0] I_10_2,
  input  [15:0] I_11_0,
  input  [15:0] I_11_1,
  input  [15:0] I_11_2,
  input  [15:0] I_12_0,
  input  [15:0] I_12_1,
  input  [15:0] I_12_2,
  input  [15:0] I_13_0,
  input  [15:0] I_13_1,
  input  [15:0] I_13_2,
  input  [15:0] I_14_0,
  input  [15:0] I_14_1,
  input  [15:0] I_14_2,
  input  [15:0] I_15_0,
  input  [15:0] I_15_1,
  input  [15:0] I_15_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2 = I_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_3_0_2 = I_3_2; // @[Partition.scala 15:39]
  assign O_4_0_0 = I_4_0; // @[Partition.scala 15:39]
  assign O_4_0_1 = I_4_1; // @[Partition.scala 15:39]
  assign O_4_0_2 = I_4_2; // @[Partition.scala 15:39]
  assign O_5_0_0 = I_5_0; // @[Partition.scala 15:39]
  assign O_5_0_1 = I_5_1; // @[Partition.scala 15:39]
  assign O_5_0_2 = I_5_2; // @[Partition.scala 15:39]
  assign O_6_0_0 = I_6_0; // @[Partition.scala 15:39]
  assign O_6_0_1 = I_6_1; // @[Partition.scala 15:39]
  assign O_6_0_2 = I_6_2; // @[Partition.scala 15:39]
  assign O_7_0_0 = I_7_0; // @[Partition.scala 15:39]
  assign O_7_0_1 = I_7_1; // @[Partition.scala 15:39]
  assign O_7_0_2 = I_7_2; // @[Partition.scala 15:39]
  assign O_8_0_0 = I_8_0; // @[Partition.scala 15:39]
  assign O_8_0_1 = I_8_1; // @[Partition.scala 15:39]
  assign O_8_0_2 = I_8_2; // @[Partition.scala 15:39]
  assign O_9_0_0 = I_9_0; // @[Partition.scala 15:39]
  assign O_9_0_1 = I_9_1; // @[Partition.scala 15:39]
  assign O_9_0_2 = I_9_2; // @[Partition.scala 15:39]
  assign O_10_0_0 = I_10_0; // @[Partition.scala 15:39]
  assign O_10_0_1 = I_10_1; // @[Partition.scala 15:39]
  assign O_10_0_2 = I_10_2; // @[Partition.scala 15:39]
  assign O_11_0_0 = I_11_0; // @[Partition.scala 15:39]
  assign O_11_0_1 = I_11_1; // @[Partition.scala 15:39]
  assign O_11_0_2 = I_11_2; // @[Partition.scala 15:39]
  assign O_12_0_0 = I_12_0; // @[Partition.scala 15:39]
  assign O_12_0_1 = I_12_1; // @[Partition.scala 15:39]
  assign O_12_0_2 = I_12_2; // @[Partition.scala 15:39]
  assign O_13_0_0 = I_13_0; // @[Partition.scala 15:39]
  assign O_13_0_1 = I_13_1; // @[Partition.scala 15:39]
  assign O_13_0_2 = I_13_2; // @[Partition.scala 15:39]
  assign O_14_0_0 = I_14_0; // @[Partition.scala 15:39]
  assign O_14_0_1 = I_14_1; // @[Partition.scala 15:39]
  assign O_14_0_2 = I_14_2; // @[Partition.scala 15:39]
  assign O_15_0_0 = I_15_0; // @[Partition.scala 15:39]
  assign O_15_0_1 = I_15_1; // @[Partition.scala 15:39]
  assign O_15_0_2 = I_15_2; // @[Partition.scala 15:39]
endmodule
module MapT(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  input  [15:0] I_4_0,
  input  [15:0] I_4_1,
  input  [15:0] I_4_2,
  input  [15:0] I_5_0,
  input  [15:0] I_5_1,
  input  [15:0] I_5_2,
  input  [15:0] I_6_0,
  input  [15:0] I_6_1,
  input  [15:0] I_6_2,
  input  [15:0] I_7_0,
  input  [15:0] I_7_1,
  input  [15:0] I_7_2,
  input  [15:0] I_8_0,
  input  [15:0] I_8_1,
  input  [15:0] I_8_2,
  input  [15:0] I_9_0,
  input  [15:0] I_9_1,
  input  [15:0] I_9_2,
  input  [15:0] I_10_0,
  input  [15:0] I_10_1,
  input  [15:0] I_10_2,
  input  [15:0] I_11_0,
  input  [15:0] I_11_1,
  input  [15:0] I_11_2,
  input  [15:0] I_12_0,
  input  [15:0] I_12_1,
  input  [15:0] I_12_2,
  input  [15:0] I_13_0,
  input  [15:0] I_13_1,
  input  [15:0] I_13_2,
  input  [15:0] I_14_0,
  input  [15:0] I_14_1,
  input  [15:0] I_14_2,
  input  [15:0] I_15_0,
  input  [15:0] I_15_1,
  input  [15:0] I_15_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_2; // @[MapT.scala 8:20]
  PartitionS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_1_2(op_I_1_2),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_2_2(op_I_2_2),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .I_3_2(op_I_3_2),
    .I_4_0(op_I_4_0),
    .I_4_1(op_I_4_1),
    .I_4_2(op_I_4_2),
    .I_5_0(op_I_5_0),
    .I_5_1(op_I_5_1),
    .I_5_2(op_I_5_2),
    .I_6_0(op_I_6_0),
    .I_6_1(op_I_6_1),
    .I_6_2(op_I_6_2),
    .I_7_0(op_I_7_0),
    .I_7_1(op_I_7_1),
    .I_7_2(op_I_7_2),
    .I_8_0(op_I_8_0),
    .I_8_1(op_I_8_1),
    .I_8_2(op_I_8_2),
    .I_9_0(op_I_9_0),
    .I_9_1(op_I_9_1),
    .I_9_2(op_I_9_2),
    .I_10_0(op_I_10_0),
    .I_10_1(op_I_10_1),
    .I_10_2(op_I_10_2),
    .I_11_0(op_I_11_0),
    .I_11_1(op_I_11_1),
    .I_11_2(op_I_11_2),
    .I_12_0(op_I_12_0),
    .I_12_1(op_I_12_1),
    .I_12_2(op_I_12_2),
    .I_13_0(op_I_13_0),
    .I_13_1(op_I_13_1),
    .I_13_2(op_I_13_2),
    .I_14_0(op_I_14_0),
    .I_14_1(op_I_14_1),
    .I_14_2(op_I_14_2),
    .I_15_0(op_I_15_0),
    .I_15_1(op_I_15_1),
    .I_15_2(op_I_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_1_2 = I_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2 = I_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
  assign op_I_3_2 = I_3_2; // @[MapT.scala 14:10]
  assign op_I_4_0 = I_4_0; // @[MapT.scala 14:10]
  assign op_I_4_1 = I_4_1; // @[MapT.scala 14:10]
  assign op_I_4_2 = I_4_2; // @[MapT.scala 14:10]
  assign op_I_5_0 = I_5_0; // @[MapT.scala 14:10]
  assign op_I_5_1 = I_5_1; // @[MapT.scala 14:10]
  assign op_I_5_2 = I_5_2; // @[MapT.scala 14:10]
  assign op_I_6_0 = I_6_0; // @[MapT.scala 14:10]
  assign op_I_6_1 = I_6_1; // @[MapT.scala 14:10]
  assign op_I_6_2 = I_6_2; // @[MapT.scala 14:10]
  assign op_I_7_0 = I_7_0; // @[MapT.scala 14:10]
  assign op_I_7_1 = I_7_1; // @[MapT.scala 14:10]
  assign op_I_7_2 = I_7_2; // @[MapT.scala 14:10]
  assign op_I_8_0 = I_8_0; // @[MapT.scala 14:10]
  assign op_I_8_1 = I_8_1; // @[MapT.scala 14:10]
  assign op_I_8_2 = I_8_2; // @[MapT.scala 14:10]
  assign op_I_9_0 = I_9_0; // @[MapT.scala 14:10]
  assign op_I_9_1 = I_9_1; // @[MapT.scala 14:10]
  assign op_I_9_2 = I_9_2; // @[MapT.scala 14:10]
  assign op_I_10_0 = I_10_0; // @[MapT.scala 14:10]
  assign op_I_10_1 = I_10_1; // @[MapT.scala 14:10]
  assign op_I_10_2 = I_10_2; // @[MapT.scala 14:10]
  assign op_I_11_0 = I_11_0; // @[MapT.scala 14:10]
  assign op_I_11_1 = I_11_1; // @[MapT.scala 14:10]
  assign op_I_11_2 = I_11_2; // @[MapT.scala 14:10]
  assign op_I_12_0 = I_12_0; // @[MapT.scala 14:10]
  assign op_I_12_1 = I_12_1; // @[MapT.scala 14:10]
  assign op_I_12_2 = I_12_2; // @[MapT.scala 14:10]
  assign op_I_13_0 = I_13_0; // @[MapT.scala 14:10]
  assign op_I_13_1 = I_13_1; // @[MapT.scala 14:10]
  assign op_I_13_2 = I_13_2; // @[MapT.scala 14:10]
  assign op_I_14_0 = I_14_0; // @[MapT.scala 14:10]
  assign op_I_14_1 = I_14_1; // @[MapT.scala 14:10]
  assign op_I_14_2 = I_14_2; // @[MapT.scala 14:10]
  assign op_I_15_0 = I_15_0; // @[MapT.scala 14:10]
  assign op_I_15_1 = I_15_1; // @[MapT.scala 14:10]
  assign op_I_15_2 = I_15_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_8_0_0,
  input  [15:0] I_8_0_1,
  input  [15:0] I_8_0_2,
  input  [15:0] I_9_0_0,
  input  [15:0] I_9_0_1,
  input  [15:0] I_9_0_2,
  input  [15:0] I_10_0_0,
  input  [15:0] I_10_0_1,
  input  [15:0] I_10_0_2,
  input  [15:0] I_11_0_0,
  input  [15:0] I_11_0_1,
  input  [15:0] I_11_0_2,
  input  [15:0] I_12_0_0,
  input  [15:0] I_12_0_1,
  input  [15:0] I_12_0_2,
  input  [15:0] I_13_0_0,
  input  [15:0] I_13_0_1,
  input  [15:0] I_13_0_2,
  input  [15:0] I_14_0_0,
  input  [15:0] I_14_0_1,
  input  [15:0] I_14_0_2,
  input  [15:0] I_15_0_0,
  input  [15:0] I_15_0_1,
  input  [15:0] I_15_0_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_8_2,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_9_2,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_10_2,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_11_2,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_12_2,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_13_2,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_14_2,
  output [15:0] O_15_0,
  output [15:0] O_15_1,
  output [15:0] O_15_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  Remove1S other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  Remove1S other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  Remove1S other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  Remove1S other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  Remove1S other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  Remove1S other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  Remove1S other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  Remove1S other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  Remove1S other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  Remove1S other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  Remove1S other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  Remove1S other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  Remove1S other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  Remove1S other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_3_2 = other_ops_2_O_2; // @[MapS.scala 21:12]
  assign O_4_0 = other_ops_3_O_0; // @[MapS.scala 21:12]
  assign O_4_1 = other_ops_3_O_1; // @[MapS.scala 21:12]
  assign O_4_2 = other_ops_3_O_2; // @[MapS.scala 21:12]
  assign O_5_0 = other_ops_4_O_0; // @[MapS.scala 21:12]
  assign O_5_1 = other_ops_4_O_1; // @[MapS.scala 21:12]
  assign O_5_2 = other_ops_4_O_2; // @[MapS.scala 21:12]
  assign O_6_0 = other_ops_5_O_0; // @[MapS.scala 21:12]
  assign O_6_1 = other_ops_5_O_1; // @[MapS.scala 21:12]
  assign O_6_2 = other_ops_5_O_2; // @[MapS.scala 21:12]
  assign O_7_0 = other_ops_6_O_0; // @[MapS.scala 21:12]
  assign O_7_1 = other_ops_6_O_1; // @[MapS.scala 21:12]
  assign O_7_2 = other_ops_6_O_2; // @[MapS.scala 21:12]
  assign O_8_0 = other_ops_7_O_0; // @[MapS.scala 21:12]
  assign O_8_1 = other_ops_7_O_1; // @[MapS.scala 21:12]
  assign O_8_2 = other_ops_7_O_2; // @[MapS.scala 21:12]
  assign O_9_0 = other_ops_8_O_0; // @[MapS.scala 21:12]
  assign O_9_1 = other_ops_8_O_1; // @[MapS.scala 21:12]
  assign O_9_2 = other_ops_8_O_2; // @[MapS.scala 21:12]
  assign O_10_0 = other_ops_9_O_0; // @[MapS.scala 21:12]
  assign O_10_1 = other_ops_9_O_1; // @[MapS.scala 21:12]
  assign O_10_2 = other_ops_9_O_2; // @[MapS.scala 21:12]
  assign O_11_0 = other_ops_10_O_0; // @[MapS.scala 21:12]
  assign O_11_1 = other_ops_10_O_1; // @[MapS.scala 21:12]
  assign O_11_2 = other_ops_10_O_2; // @[MapS.scala 21:12]
  assign O_12_0 = other_ops_11_O_0; // @[MapS.scala 21:12]
  assign O_12_1 = other_ops_11_O_1; // @[MapS.scala 21:12]
  assign O_12_2 = other_ops_11_O_2; // @[MapS.scala 21:12]
  assign O_13_0 = other_ops_12_O_0; // @[MapS.scala 21:12]
  assign O_13_1 = other_ops_12_O_1; // @[MapS.scala 21:12]
  assign O_13_2 = other_ops_12_O_2; // @[MapS.scala 21:12]
  assign O_14_0 = other_ops_13_O_0; // @[MapS.scala 21:12]
  assign O_14_1 = other_ops_13_O_1; // @[MapS.scala 21:12]
  assign O_14_2 = other_ops_13_O_2; // @[MapS.scala 21:12]
  assign O_15_0 = other_ops_14_O_0; // @[MapS.scala 21:12]
  assign O_15_1 = other_ops_14_O_1; // @[MapS.scala 21:12]
  assign O_15_2 = other_ops_14_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
endmodule
module MapT_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_8_0_0,
  input  [15:0] I_8_0_1,
  input  [15:0] I_8_0_2,
  input  [15:0] I_9_0_0,
  input  [15:0] I_9_0_1,
  input  [15:0] I_9_0_2,
  input  [15:0] I_10_0_0,
  input  [15:0] I_10_0_1,
  input  [15:0] I_10_0_2,
  input  [15:0] I_11_0_0,
  input  [15:0] I_11_0_1,
  input  [15:0] I_11_0_2,
  input  [15:0] I_12_0_0,
  input  [15:0] I_12_0_1,
  input  [15:0] I_12_0_2,
  input  [15:0] I_13_0_0,
  input  [15:0] I_13_0_1,
  input  [15:0] I_13_0_2,
  input  [15:0] I_14_0_0,
  input  [15:0] I_14_0_1,
  input  [15:0] I_14_0_2,
  input  [15:0] I_15_0_0,
  input  [15:0] I_15_0_1,
  input  [15:0] I_15_0_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_8_2,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_9_2,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_10_2,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_11_2,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_12_2,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_13_2,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_14_2,
  output [15:0] O_15_0,
  output [15:0] O_15_1,
  output [15:0] O_15_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_2; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_8_2(op_O_8_2),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_9_2(op_O_9_2),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_10_2(op_O_10_2),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_11_2(op_O_11_2),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_12_2(op_O_12_2),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_13_2(op_O_13_2),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_14_2(op_O_14_2),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1),
    .O_15_2(op_O_15_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_0_2 = op_O_0_2; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_1_2 = op_O_1_2; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_2_2 = op_O_2_2; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign O_3_2 = op_O_3_2; // @[MapT.scala 15:7]
  assign O_4_0 = op_O_4_0; // @[MapT.scala 15:7]
  assign O_4_1 = op_O_4_1; // @[MapT.scala 15:7]
  assign O_4_2 = op_O_4_2; // @[MapT.scala 15:7]
  assign O_5_0 = op_O_5_0; // @[MapT.scala 15:7]
  assign O_5_1 = op_O_5_1; // @[MapT.scala 15:7]
  assign O_5_2 = op_O_5_2; // @[MapT.scala 15:7]
  assign O_6_0 = op_O_6_0; // @[MapT.scala 15:7]
  assign O_6_1 = op_O_6_1; // @[MapT.scala 15:7]
  assign O_6_2 = op_O_6_2; // @[MapT.scala 15:7]
  assign O_7_0 = op_O_7_0; // @[MapT.scala 15:7]
  assign O_7_1 = op_O_7_1; // @[MapT.scala 15:7]
  assign O_7_2 = op_O_7_2; // @[MapT.scala 15:7]
  assign O_8_0 = op_O_8_0; // @[MapT.scala 15:7]
  assign O_8_1 = op_O_8_1; // @[MapT.scala 15:7]
  assign O_8_2 = op_O_8_2; // @[MapT.scala 15:7]
  assign O_9_0 = op_O_9_0; // @[MapT.scala 15:7]
  assign O_9_1 = op_O_9_1; // @[MapT.scala 15:7]
  assign O_9_2 = op_O_9_2; // @[MapT.scala 15:7]
  assign O_10_0 = op_O_10_0; // @[MapT.scala 15:7]
  assign O_10_1 = op_O_10_1; // @[MapT.scala 15:7]
  assign O_10_2 = op_O_10_2; // @[MapT.scala 15:7]
  assign O_11_0 = op_O_11_0; // @[MapT.scala 15:7]
  assign O_11_1 = op_O_11_1; // @[MapT.scala 15:7]
  assign O_11_2 = op_O_11_2; // @[MapT.scala 15:7]
  assign O_12_0 = op_O_12_0; // @[MapT.scala 15:7]
  assign O_12_1 = op_O_12_1; // @[MapT.scala 15:7]
  assign O_12_2 = op_O_12_2; // @[MapT.scala 15:7]
  assign O_13_0 = op_O_13_0; // @[MapT.scala 15:7]
  assign O_13_1 = op_O_13_1; // @[MapT.scala 15:7]
  assign O_13_2 = op_O_13_2; // @[MapT.scala 15:7]
  assign O_14_0 = op_O_14_0; // @[MapT.scala 15:7]
  assign O_14_1 = op_O_14_1; // @[MapT.scala 15:7]
  assign O_14_2 = op_O_14_2; // @[MapT.scala 15:7]
  assign O_15_0 = op_O_15_0; // @[MapT.scala 15:7]
  assign O_15_1 = op_O_15_1; // @[MapT.scala 15:7]
  assign O_15_2 = op_O_15_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
endmodule
module FIFO_5(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  input  [15:0] I_4_0,
  input  [15:0] I_4_1,
  input  [15:0] I_4_2,
  input  [15:0] I_5_0,
  input  [15:0] I_5_1,
  input  [15:0] I_5_2,
  input  [15:0] I_6_0,
  input  [15:0] I_6_1,
  input  [15:0] I_6_2,
  input  [15:0] I_7_0,
  input  [15:0] I_7_1,
  input  [15:0] I_7_2,
  input  [15:0] I_8_0,
  input  [15:0] I_8_1,
  input  [15:0] I_8_2,
  input  [15:0] I_9_0,
  input  [15:0] I_9_1,
  input  [15:0] I_9_2,
  input  [15:0] I_10_0,
  input  [15:0] I_10_1,
  input  [15:0] I_10_2,
  input  [15:0] I_11_0,
  input  [15:0] I_11_1,
  input  [15:0] I_11_2,
  input  [15:0] I_12_0,
  input  [15:0] I_12_1,
  input  [15:0] I_12_2,
  input  [15:0] I_13_0,
  input  [15:0] I_13_1,
  input  [15:0] I_13_2,
  input  [15:0] I_14_0,
  input  [15:0] I_14_1,
  input  [15:0] I_14_2,
  input  [15:0] I_15_0,
  input  [15:0] I_15_1,
  input  [15:0] I_15_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_8_2,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_9_2,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_10_2,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_11_2,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_12_2,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_13_2,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_14_2,
  output [15:0] O_15_0,
  output [15:0] O_15_1,
  output [15:0] O_15_2
);
  reg [15:0] _T__0_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [15:0] _T__0_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [15:0] _T__0_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [15:0] _T__1_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [15:0] _T__1_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [15:0] _T__1_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [15:0] _T__2_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [15:0] _T__2_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [15:0] _T__2_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [15:0] _T__3_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [15:0] _T__3_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [15:0] _T__3_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [15:0] _T__4_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [15:0] _T__4_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [15:0] _T__4_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [15:0] _T__5_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg [15:0] _T__5_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_16;
  reg [15:0] _T__5_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_17;
  reg [15:0] _T__6_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_18;
  reg [15:0] _T__6_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_19;
  reg [15:0] _T__6_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_20;
  reg [15:0] _T__7_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_21;
  reg [15:0] _T__7_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_22;
  reg [15:0] _T__7_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_23;
  reg [15:0] _T__8_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_24;
  reg [15:0] _T__8_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_25;
  reg [15:0] _T__8_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_26;
  reg [15:0] _T__9_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_27;
  reg [15:0] _T__9_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_28;
  reg [15:0] _T__9_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_29;
  reg [15:0] _T__10_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_30;
  reg [15:0] _T__10_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_31;
  reg [15:0] _T__10_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_32;
  reg [15:0] _T__11_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_33;
  reg [15:0] _T__11_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_34;
  reg [15:0] _T__11_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_35;
  reg [15:0] _T__12_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_36;
  reg [15:0] _T__12_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_37;
  reg [15:0] _T__12_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_38;
  reg [15:0] _T__13_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_39;
  reg [15:0] _T__13_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_40;
  reg [15:0] _T__13_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_41;
  reg [15:0] _T__14_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_42;
  reg [15:0] _T__14_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_43;
  reg [15:0] _T__14_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_44;
  reg [15:0] _T__15_0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_45;
  reg [15:0] _T__15_1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_46;
  reg [15:0] _T__15_2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_47;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_48;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0_0 = _T__0_0; // @[FIFO.scala 14:7]
  assign O_0_1 = _T__0_1; // @[FIFO.scala 14:7]
  assign O_0_2 = _T__0_2; // @[FIFO.scala 14:7]
  assign O_1_0 = _T__1_0; // @[FIFO.scala 14:7]
  assign O_1_1 = _T__1_1; // @[FIFO.scala 14:7]
  assign O_1_2 = _T__1_2; // @[FIFO.scala 14:7]
  assign O_2_0 = _T__2_0; // @[FIFO.scala 14:7]
  assign O_2_1 = _T__2_1; // @[FIFO.scala 14:7]
  assign O_2_2 = _T__2_2; // @[FIFO.scala 14:7]
  assign O_3_0 = _T__3_0; // @[FIFO.scala 14:7]
  assign O_3_1 = _T__3_1; // @[FIFO.scala 14:7]
  assign O_3_2 = _T__3_2; // @[FIFO.scala 14:7]
  assign O_4_0 = _T__4_0; // @[FIFO.scala 14:7]
  assign O_4_1 = _T__4_1; // @[FIFO.scala 14:7]
  assign O_4_2 = _T__4_2; // @[FIFO.scala 14:7]
  assign O_5_0 = _T__5_0; // @[FIFO.scala 14:7]
  assign O_5_1 = _T__5_1; // @[FIFO.scala 14:7]
  assign O_5_2 = _T__5_2; // @[FIFO.scala 14:7]
  assign O_6_0 = _T__6_0; // @[FIFO.scala 14:7]
  assign O_6_1 = _T__6_1; // @[FIFO.scala 14:7]
  assign O_6_2 = _T__6_2; // @[FIFO.scala 14:7]
  assign O_7_0 = _T__7_0; // @[FIFO.scala 14:7]
  assign O_7_1 = _T__7_1; // @[FIFO.scala 14:7]
  assign O_7_2 = _T__7_2; // @[FIFO.scala 14:7]
  assign O_8_0 = _T__8_0; // @[FIFO.scala 14:7]
  assign O_8_1 = _T__8_1; // @[FIFO.scala 14:7]
  assign O_8_2 = _T__8_2; // @[FIFO.scala 14:7]
  assign O_9_0 = _T__9_0; // @[FIFO.scala 14:7]
  assign O_9_1 = _T__9_1; // @[FIFO.scala 14:7]
  assign O_9_2 = _T__9_2; // @[FIFO.scala 14:7]
  assign O_10_0 = _T__10_0; // @[FIFO.scala 14:7]
  assign O_10_1 = _T__10_1; // @[FIFO.scala 14:7]
  assign O_10_2 = _T__10_2; // @[FIFO.scala 14:7]
  assign O_11_0 = _T__11_0; // @[FIFO.scala 14:7]
  assign O_11_1 = _T__11_1; // @[FIFO.scala 14:7]
  assign O_11_2 = _T__11_2; // @[FIFO.scala 14:7]
  assign O_12_0 = _T__12_0; // @[FIFO.scala 14:7]
  assign O_12_1 = _T__12_1; // @[FIFO.scala 14:7]
  assign O_12_2 = _T__12_2; // @[FIFO.scala 14:7]
  assign O_13_0 = _T__13_0; // @[FIFO.scala 14:7]
  assign O_13_1 = _T__13_1; // @[FIFO.scala 14:7]
  assign O_13_2 = _T__13_2; // @[FIFO.scala 14:7]
  assign O_14_0 = _T__14_0; // @[FIFO.scala 14:7]
  assign O_14_1 = _T__14_1; // @[FIFO.scala 14:7]
  assign O_14_2 = _T__14_2; // @[FIFO.scala 14:7]
  assign O_15_0 = _T__15_0; // @[FIFO.scala 14:7]
  assign O_15_1 = _T__15_1; // @[FIFO.scala 14:7]
  assign O_15_2 = _T__15_2; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__0_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__1_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__1_1 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__1_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__2_0 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__2_1 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__2_2 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__3_0 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__3_1 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__3_2 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__4_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__4_1 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__4_2 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__5_0 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T__5_1 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T__5_2 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__6_0 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__6_1 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T__6_2 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T__7_0 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__7_1 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__7_2 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T__8_0 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T__8_1 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__8_2 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__9_0 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T__9_1 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T__9_2 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__10_0 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__10_1 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T__10_2 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T__11_0 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__11_1 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__11_2 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T__12_0 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T__12_1 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__12_2 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__13_0 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T__13_1 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T__13_2 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T__14_0 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T__14_1 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T__14_2 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T__15_0 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T__15_1 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T__15_2 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0_0 <= I_0_0;
    _T__0_1 <= I_0_1;
    _T__0_2 <= I_0_2;
    _T__1_0 <= I_1_0;
    _T__1_1 <= I_1_1;
    _T__1_2 <= I_1_2;
    _T__2_0 <= I_2_0;
    _T__2_1 <= I_2_1;
    _T__2_2 <= I_2_2;
    _T__3_0 <= I_3_0;
    _T__3_1 <= I_3_1;
    _T__3_2 <= I_3_2;
    _T__4_0 <= I_4_0;
    _T__4_1 <= I_4_1;
    _T__4_2 <= I_4_2;
    _T__5_0 <= I_5_0;
    _T__5_1 <= I_5_1;
    _T__5_2 <= I_5_2;
    _T__6_0 <= I_6_0;
    _T__6_1 <= I_6_1;
    _T__6_2 <= I_6_2;
    _T__7_0 <= I_7_0;
    _T__7_1 <= I_7_1;
    _T__7_2 <= I_7_2;
    _T__8_0 <= I_8_0;
    _T__8_1 <= I_8_1;
    _T__8_2 <= I_8_2;
    _T__9_0 <= I_9_0;
    _T__9_1 <= I_9_1;
    _T__9_2 <= I_9_2;
    _T__10_0 <= I_10_0;
    _T__10_1 <= I_10_1;
    _T__10_2 <= I_10_2;
    _T__11_0 <= I_11_0;
    _T__11_1 <= I_11_1;
    _T__11_2 <= I_11_2;
    _T__12_0 <= I_12_0;
    _T__12_1 <= I_12_1;
    _T__12_2 <= I_12_2;
    _T__13_0 <= I_13_0;
    _T__13_1 <= I_13_1;
    _T__13_2 <= I_13_2;
    _T__14_0 <= I_14_0;
    _T__14_1 <= I_14_1;
    _T__14_2 <= I_14_2;
    _T__15_0 <= I_15_0;
    _T__15_1 <= I_15_1;
    _T__15_2 <= I_15_2;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module SSeqTupleCreator_2(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_3_2,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_4_2,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_5_2,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_6_2,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I0_7_2,
  input  [15:0] I0_8_0,
  input  [15:0] I0_8_1,
  input  [15:0] I0_8_2,
  input  [15:0] I0_9_0,
  input  [15:0] I0_9_1,
  input  [15:0] I0_9_2,
  input  [15:0] I0_10_0,
  input  [15:0] I0_10_1,
  input  [15:0] I0_10_2,
  input  [15:0] I0_11_0,
  input  [15:0] I0_11_1,
  input  [15:0] I0_11_2,
  input  [15:0] I0_12_0,
  input  [15:0] I0_12_1,
  input  [15:0] I0_12_2,
  input  [15:0] I0_13_0,
  input  [15:0] I0_13_1,
  input  [15:0] I0_13_2,
  input  [15:0] I0_14_0,
  input  [15:0] I0_14_1,
  input  [15:0] I0_14_2,
  input  [15:0] I0_15_0,
  input  [15:0] I0_15_1,
  input  [15:0] I0_15_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  input  [15:0] I1_8_0,
  input  [15:0] I1_8_1,
  input  [15:0] I1_8_2,
  input  [15:0] I1_9_0,
  input  [15:0] I1_9_1,
  input  [15:0] I1_9_2,
  input  [15:0] I1_10_0,
  input  [15:0] I1_10_1,
  input  [15:0] I1_10_2,
  input  [15:0] I1_11_0,
  input  [15:0] I1_11_1,
  input  [15:0] I1_11_2,
  input  [15:0] I1_12_0,
  input  [15:0] I1_12_1,
  input  [15:0] I1_12_2,
  input  [15:0] I1_13_0,
  input  [15:0] I1_13_1,
  input  [15:0] I1_13_2,
  input  [15:0] I1_14_0,
  input  [15:0] I1_14_1,
  input  [15:0] I1_14_2,
  input  [15:0] I1_15_0,
  input  [15:0] I1_15_1,
  input  [15:0] I1_15_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_8_1_0,
  output [15:0] O_8_1_1,
  output [15:0] O_8_1_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_9_1_0,
  output [15:0] O_9_1_1,
  output [15:0] O_9_1_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_10_1_0,
  output [15:0] O_10_1_1,
  output [15:0] O_10_1_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_11_1_0,
  output [15:0] O_11_1_1,
  output [15:0] O_11_1_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_12_1_0,
  output [15:0] O_12_1_1,
  output [15:0] O_12_1_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_13_1_0,
  output [15:0] O_13_1_1,
  output [15:0] O_13_1_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_14_1_0,
  output [15:0] O_14_1_1,
  output [15:0] O_14_1_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2,
  output [15:0] O_15_1_0,
  output [15:0] O_15_1_1,
  output [15:0] O_15_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I0_2(other_ops_2_I0_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I0_2(other_ops_3_I0_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I0_2(other_ops_4_I0_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I0_2(other_ops_5_I0_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I0_2(other_ops_6_I0_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I0_2(other_ops_7_I0_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I0_2(other_ops_8_I0_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I0_2(other_ops_9_I0_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I0_2(other_ops_10_I0_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I0_2(other_ops_11_I0_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I0_2(other_ops_12_I0_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I0_2(other_ops_13_I0_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I0_2(other_ops_14_I0_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2 = I0_3_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2 = I0_4_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2 = I0_5_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2 = I0_6_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2 = I0_7_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_2 = I0_8_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_2 = I0_9_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_2 = I0_10_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_2 = I0_11_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_2 = I0_12_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_2 = I0_13_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_2 = I0_14_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_2 = I0_15_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  input  [15:0] I0_3_0,
  input  [15:0] I0_3_1,
  input  [15:0] I0_3_2,
  input  [15:0] I0_4_0,
  input  [15:0] I0_4_1,
  input  [15:0] I0_4_2,
  input  [15:0] I0_5_0,
  input  [15:0] I0_5_1,
  input  [15:0] I0_5_2,
  input  [15:0] I0_6_0,
  input  [15:0] I0_6_1,
  input  [15:0] I0_6_2,
  input  [15:0] I0_7_0,
  input  [15:0] I0_7_1,
  input  [15:0] I0_7_2,
  input  [15:0] I0_8_0,
  input  [15:0] I0_8_1,
  input  [15:0] I0_8_2,
  input  [15:0] I0_9_0,
  input  [15:0] I0_9_1,
  input  [15:0] I0_9_2,
  input  [15:0] I0_10_0,
  input  [15:0] I0_10_1,
  input  [15:0] I0_10_2,
  input  [15:0] I0_11_0,
  input  [15:0] I0_11_1,
  input  [15:0] I0_11_2,
  input  [15:0] I0_12_0,
  input  [15:0] I0_12_1,
  input  [15:0] I0_12_2,
  input  [15:0] I0_13_0,
  input  [15:0] I0_13_1,
  input  [15:0] I0_13_2,
  input  [15:0] I0_14_0,
  input  [15:0] I0_14_1,
  input  [15:0] I0_14_2,
  input  [15:0] I0_15_0,
  input  [15:0] I0_15_1,
  input  [15:0] I0_15_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  input  [15:0] I1_8_0,
  input  [15:0] I1_8_1,
  input  [15:0] I1_8_2,
  input  [15:0] I1_9_0,
  input  [15:0] I1_9_1,
  input  [15:0] I1_9_2,
  input  [15:0] I1_10_0,
  input  [15:0] I1_10_1,
  input  [15:0] I1_10_2,
  input  [15:0] I1_11_0,
  input  [15:0] I1_11_1,
  input  [15:0] I1_11_2,
  input  [15:0] I1_12_0,
  input  [15:0] I1_12_1,
  input  [15:0] I1_12_2,
  input  [15:0] I1_13_0,
  input  [15:0] I1_13_1,
  input  [15:0] I1_13_2,
  input  [15:0] I1_14_0,
  input  [15:0] I1_14_1,
  input  [15:0] I1_14_2,
  input  [15:0] I1_15_0,
  input  [15:0] I1_15_1,
  input  [15:0] I1_15_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_8_1_0,
  output [15:0] O_8_1_1,
  output [15:0] O_8_1_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_9_1_0,
  output [15:0] O_9_1_1,
  output [15:0] O_9_1_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_10_1_0,
  output [15:0] O_10_1_1,
  output [15:0] O_10_1_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_11_1_0,
  output [15:0] O_11_1_1,
  output [15:0] O_11_1_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_12_1_0,
  output [15:0] O_12_1_1,
  output [15:0] O_12_1_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_13_1_0,
  output [15:0] O_13_1_1,
  output [15:0] O_13_1_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_14_1_0,
  output [15:0] O_14_1_1,
  output [15:0] O_14_1_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2,
  output [15:0] O_15_1_0,
  output [15:0] O_15_1_1,
  output [15:0] O_15_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1_2; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_0_2(op_I0_0_2),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_1_2(op_I0_1_2),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_2_2(op_I0_2_2),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_3_2(op_I0_3_2),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_4_2(op_I0_4_2),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_5_2(op_I0_5_2),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_6_2(op_I0_6_2),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_7_2(op_I0_7_2),
    .I0_8_0(op_I0_8_0),
    .I0_8_1(op_I0_8_1),
    .I0_8_2(op_I0_8_2),
    .I0_9_0(op_I0_9_0),
    .I0_9_1(op_I0_9_1),
    .I0_9_2(op_I0_9_2),
    .I0_10_0(op_I0_10_0),
    .I0_10_1(op_I0_10_1),
    .I0_10_2(op_I0_10_2),
    .I0_11_0(op_I0_11_0),
    .I0_11_1(op_I0_11_1),
    .I0_11_2(op_I0_11_2),
    .I0_12_0(op_I0_12_0),
    .I0_12_1(op_I0_12_1),
    .I0_12_2(op_I0_12_2),
    .I0_13_0(op_I0_13_0),
    .I0_13_1(op_I0_13_1),
    .I0_13_2(op_I0_13_2),
    .I0_14_0(op_I0_14_0),
    .I0_14_1(op_I0_14_1),
    .I0_14_2(op_I0_14_2),
    .I0_15_0(op_I0_15_0),
    .I0_15_1(op_I0_15_1),
    .I0_15_2(op_I0_15_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .I1_8_0(op_I1_8_0),
    .I1_8_1(op_I1_8_1),
    .I1_8_2(op_I1_8_2),
    .I1_9_0(op_I1_9_0),
    .I1_9_1(op_I1_9_1),
    .I1_9_2(op_I1_9_2),
    .I1_10_0(op_I1_10_0),
    .I1_10_1(op_I1_10_1),
    .I1_10_2(op_I1_10_2),
    .I1_11_0(op_I1_11_0),
    .I1_11_1(op_I1_11_1),
    .I1_11_2(op_I1_11_2),
    .I1_12_0(op_I1_12_0),
    .I1_12_1(op_I1_12_1),
    .I1_12_2(op_I1_12_2),
    .I1_13_0(op_I1_13_0),
    .I1_13_1(op_I1_13_1),
    .I1_13_2(op_I1_13_2),
    .I1_14_0(op_I1_14_0),
    .I1_14_1(op_I1_14_1),
    .I1_14_2(op_I1_14_2),
    .I1_15_0(op_I1_15_0),
    .I1_15_1(op_I1_15_1),
    .I1_15_2(op_I1_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_1 = op_O_8_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_2 = op_O_8_0_2; // @[Map2T.scala 17:7]
  assign O_8_1_0 = op_O_8_1_0; // @[Map2T.scala 17:7]
  assign O_8_1_1 = op_O_8_1_1; // @[Map2T.scala 17:7]
  assign O_8_1_2 = op_O_8_1_2; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_1 = op_O_9_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_2 = op_O_9_0_2; // @[Map2T.scala 17:7]
  assign O_9_1_0 = op_O_9_1_0; // @[Map2T.scala 17:7]
  assign O_9_1_1 = op_O_9_1_1; // @[Map2T.scala 17:7]
  assign O_9_1_2 = op_O_9_1_2; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_1 = op_O_10_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_2 = op_O_10_0_2; // @[Map2T.scala 17:7]
  assign O_10_1_0 = op_O_10_1_0; // @[Map2T.scala 17:7]
  assign O_10_1_1 = op_O_10_1_1; // @[Map2T.scala 17:7]
  assign O_10_1_2 = op_O_10_1_2; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_1 = op_O_11_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_2 = op_O_11_0_2; // @[Map2T.scala 17:7]
  assign O_11_1_0 = op_O_11_1_0; // @[Map2T.scala 17:7]
  assign O_11_1_1 = op_O_11_1_1; // @[Map2T.scala 17:7]
  assign O_11_1_2 = op_O_11_1_2; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_1 = op_O_12_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_2 = op_O_12_0_2; // @[Map2T.scala 17:7]
  assign O_12_1_0 = op_O_12_1_0; // @[Map2T.scala 17:7]
  assign O_12_1_1 = op_O_12_1_1; // @[Map2T.scala 17:7]
  assign O_12_1_2 = op_O_12_1_2; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_1 = op_O_13_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_2 = op_O_13_0_2; // @[Map2T.scala 17:7]
  assign O_13_1_0 = op_O_13_1_0; // @[Map2T.scala 17:7]
  assign O_13_1_1 = op_O_13_1_1; // @[Map2T.scala 17:7]
  assign O_13_1_2 = op_O_13_1_2; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_1 = op_O_14_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_2 = op_O_14_0_2; // @[Map2T.scala 17:7]
  assign O_14_1_0 = op_O_14_1_0; // @[Map2T.scala 17:7]
  assign O_14_1_1 = op_O_14_1_1; // @[Map2T.scala 17:7]
  assign O_14_1_2 = op_O_14_1_2; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_1 = op_O_15_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_2 = op_O_15_0_2; // @[Map2T.scala 17:7]
  assign O_15_1_0 = op_O_15_1_0; // @[Map2T.scala 17:7]
  assign O_15_1_1 = op_O_15_1_1; // @[Map2T.scala 17:7]
  assign O_15_1_2 = op_O_15_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2 = I0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2 = I0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2 = I0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2 = I0_3_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_4_2 = I0_4_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_5_2 = I0_5_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_6_2 = I0_6_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_7_2 = I0_7_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0 = I0_8_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1 = I0_8_1; // @[Map2T.scala 15:11]
  assign op_I0_8_2 = I0_8_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0 = I0_9_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1 = I0_9_1; // @[Map2T.scala 15:11]
  assign op_I0_9_2 = I0_9_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0 = I0_10_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1 = I0_10_1; // @[Map2T.scala 15:11]
  assign op_I0_10_2 = I0_10_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0 = I0_11_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1 = I0_11_1; // @[Map2T.scala 15:11]
  assign op_I0_11_2 = I0_11_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0 = I0_12_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1 = I0_12_1; // @[Map2T.scala 15:11]
  assign op_I0_12_2 = I0_12_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0 = I0_13_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1 = I0_13_1; // @[Map2T.scala 15:11]
  assign op_I0_13_2 = I0_13_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0 = I0_14_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1 = I0_14_1; // @[Map2T.scala 15:11]
  assign op_I0_14_2 = I0_14_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0 = I0_15_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1 = I0_15_1; // @[Map2T.scala 15:11]
  assign op_I0_15_2 = I0_15_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0 = I1_8_0; // @[Map2T.scala 16:11]
  assign op_I1_8_1 = I1_8_1; // @[Map2T.scala 16:11]
  assign op_I1_8_2 = I1_8_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0 = I1_9_0; // @[Map2T.scala 16:11]
  assign op_I1_9_1 = I1_9_1; // @[Map2T.scala 16:11]
  assign op_I1_9_2 = I1_9_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0 = I1_10_0; // @[Map2T.scala 16:11]
  assign op_I1_10_1 = I1_10_1; // @[Map2T.scala 16:11]
  assign op_I1_10_2 = I1_10_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0 = I1_11_0; // @[Map2T.scala 16:11]
  assign op_I1_11_1 = I1_11_1; // @[Map2T.scala 16:11]
  assign op_I1_11_2 = I1_11_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0 = I1_12_0; // @[Map2T.scala 16:11]
  assign op_I1_12_1 = I1_12_1; // @[Map2T.scala 16:11]
  assign op_I1_12_2 = I1_12_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0 = I1_13_0; // @[Map2T.scala 16:11]
  assign op_I1_13_1 = I1_13_1; // @[Map2T.scala 16:11]
  assign op_I1_13_2 = I1_13_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0 = I1_14_0; // @[Map2T.scala 16:11]
  assign op_I1_14_1 = I1_14_1; // @[Map2T.scala 16:11]
  assign op_I1_14_2 = I1_14_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0 = I1_15_0; // @[Map2T.scala 16:11]
  assign op_I1_15_1 = I1_15_1; // @[Map2T.scala 16:11]
  assign op_I1_15_2 = I1_15_2; // @[Map2T.scala 16:11]
endmodule
module FIFO_8(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  input  [15:0] I_3_0,
  input  [15:0] I_3_1,
  input  [15:0] I_3_2,
  input  [15:0] I_4_0,
  input  [15:0] I_4_1,
  input  [15:0] I_4_2,
  input  [15:0] I_5_0,
  input  [15:0] I_5_1,
  input  [15:0] I_5_2,
  input  [15:0] I_6_0,
  input  [15:0] I_6_1,
  input  [15:0] I_6_2,
  input  [15:0] I_7_0,
  input  [15:0] I_7_1,
  input  [15:0] I_7_2,
  input  [15:0] I_8_0,
  input  [15:0] I_8_1,
  input  [15:0] I_8_2,
  input  [15:0] I_9_0,
  input  [15:0] I_9_1,
  input  [15:0] I_9_2,
  input  [15:0] I_10_0,
  input  [15:0] I_10_1,
  input  [15:0] I_10_2,
  input  [15:0] I_11_0,
  input  [15:0] I_11_1,
  input  [15:0] I_11_2,
  input  [15:0] I_12_0,
  input  [15:0] I_12_1,
  input  [15:0] I_12_2,
  input  [15:0] I_13_0,
  input  [15:0] I_13_1,
  input  [15:0] I_13_2,
  input  [15:0] I_14_0,
  input  [15:0] I_14_1,
  input  [15:0] I_14_2,
  input  [15:0] I_15_0,
  input  [15:0] I_15_1,
  input  [15:0] I_15_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2,
  output [15:0] O_3_0,
  output [15:0] O_3_1,
  output [15:0] O_3_2,
  output [15:0] O_4_0,
  output [15:0] O_4_1,
  output [15:0] O_4_2,
  output [15:0] O_5_0,
  output [15:0] O_5_1,
  output [15:0] O_5_2,
  output [15:0] O_6_0,
  output [15:0] O_6_1,
  output [15:0] O_6_2,
  output [15:0] O_7_0,
  output [15:0] O_7_1,
  output [15:0] O_7_2,
  output [15:0] O_8_0,
  output [15:0] O_8_1,
  output [15:0] O_8_2,
  output [15:0] O_9_0,
  output [15:0] O_9_1,
  output [15:0] O_9_2,
  output [15:0] O_10_0,
  output [15:0] O_10_1,
  output [15:0] O_10_2,
  output [15:0] O_11_0,
  output [15:0] O_11_1,
  output [15:0] O_11_2,
  output [15:0] O_12_0,
  output [15:0] O_12_1,
  output [15:0] O_12_2,
  output [15:0] O_13_0,
  output [15:0] O_13_1,
  output [15:0] O_13_2,
  output [15:0] O_14_0,
  output [15:0] O_14_1,
  output [15:0] O_14_2,
  output [15:0] O_15_0,
  output [15:0] O_15_1,
  output [15:0] O_15_2
);
  reg [15:0] _T__0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [15:0] _T__0_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [15:0] _T__0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__0_0__T_17_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T__0_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [15:0] _T__0_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_4;
  wire [15:0] _T__0_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_5;
  wire [15:0] _T__0_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__0_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__0_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__0_1__T_17_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [1:0] _T__0_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [15:0] _T__0_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_8;
  wire [15:0] _T__0_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_9;
  wire [15:0] _T__0_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__0_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__0_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__0_2__T_17_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [1:0] _T__0_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [15:0] _T__1_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_12;
  wire [15:0] _T__1_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_13;
  wire [15:0] _T__1_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__1_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__1_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__1_0__T_17_en_pipe_0;
  reg [31:0] _RAND_14;
  reg [1:0] _T__1_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [15:0] _T__1_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_16;
  wire [15:0] _T__1_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_17;
  wire [15:0] _T__1_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__1_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__1_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__1_1__T_17_en_pipe_0;
  reg [31:0] _RAND_18;
  reg [1:0] _T__1_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [15:0] _T__1_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_20;
  wire [15:0] _T__1_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_21;
  wire [15:0] _T__1_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__1_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__1_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__1_2__T_17_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [1:0] _T__1_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [15:0] _T__2_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_24;
  wire [15:0] _T__2_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_25;
  wire [15:0] _T__2_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__2_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__2_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__2_0__T_17_en_pipe_0;
  reg [31:0] _RAND_26;
  reg [1:0] _T__2_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_27;
  reg [15:0] _T__2_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_28;
  wire [15:0] _T__2_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_29;
  wire [15:0] _T__2_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__2_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__2_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__2_1__T_17_en_pipe_0;
  reg [31:0] _RAND_30;
  reg [1:0] _T__2_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_31;
  reg [15:0] _T__2_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_32;
  wire [15:0] _T__2_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_33;
  wire [15:0] _T__2_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__2_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__2_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__2_2__T_17_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [1:0] _T__2_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [15:0] _T__3_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_36;
  wire [15:0] _T__3_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_37;
  wire [15:0] _T__3_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__3_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__3_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__3_0__T_17_en_pipe_0;
  reg [31:0] _RAND_38;
  reg [1:0] _T__3_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_39;
  reg [15:0] _T__3_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_40;
  wire [15:0] _T__3_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_41;
  wire [15:0] _T__3_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__3_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__3_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__3_1__T_17_en_pipe_0;
  reg [31:0] _RAND_42;
  reg [1:0] _T__3_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_43;
  reg [15:0] _T__3_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_44;
  wire [15:0] _T__3_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_45;
  wire [15:0] _T__3_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__3_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__3_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__3_2__T_17_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [1:0] _T__3_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [15:0] _T__4_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_48;
  wire [15:0] _T__4_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_49;
  wire [15:0] _T__4_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__4_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__4_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__4_0__T_17_en_pipe_0;
  reg [31:0] _RAND_50;
  reg [1:0] _T__4_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_51;
  reg [15:0] _T__4_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_52;
  wire [15:0] _T__4_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_53;
  wire [15:0] _T__4_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__4_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__4_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__4_1__T_17_en_pipe_0;
  reg [31:0] _RAND_54;
  reg [1:0] _T__4_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_55;
  reg [15:0] _T__4_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_56;
  wire [15:0] _T__4_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_57;
  wire [15:0] _T__4_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__4_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__4_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__4_2__T_17_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [1:0] _T__4_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [15:0] _T__5_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_60;
  wire [15:0] _T__5_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_61;
  wire [15:0] _T__5_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__5_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__5_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__5_0__T_17_en_pipe_0;
  reg [31:0] _RAND_62;
  reg [1:0] _T__5_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_63;
  reg [15:0] _T__5_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_64;
  wire [15:0] _T__5_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_65;
  wire [15:0] _T__5_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__5_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__5_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__5_1__T_17_en_pipe_0;
  reg [31:0] _RAND_66;
  reg [1:0] _T__5_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_67;
  reg [15:0] _T__5_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_68;
  wire [15:0] _T__5_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_69;
  wire [15:0] _T__5_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__5_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__5_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__5_2__T_17_en_pipe_0;
  reg [31:0] _RAND_70;
  reg [1:0] _T__5_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_71;
  reg [15:0] _T__6_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_72;
  wire [15:0] _T__6_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_73;
  wire [15:0] _T__6_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__6_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__6_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__6_0__T_17_en_pipe_0;
  reg [31:0] _RAND_74;
  reg [1:0] _T__6_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_75;
  reg [15:0] _T__6_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_76;
  wire [15:0] _T__6_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_77;
  wire [15:0] _T__6_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__6_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__6_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__6_1__T_17_en_pipe_0;
  reg [31:0] _RAND_78;
  reg [1:0] _T__6_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_79;
  reg [15:0] _T__6_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_80;
  wire [15:0] _T__6_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_81;
  wire [15:0] _T__6_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__6_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__6_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__6_2__T_17_en_pipe_0;
  reg [31:0] _RAND_82;
  reg [1:0] _T__6_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_83;
  reg [15:0] _T__7_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_84;
  wire [15:0] _T__7_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_85;
  wire [15:0] _T__7_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__7_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__7_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__7_0__T_17_en_pipe_0;
  reg [31:0] _RAND_86;
  reg [1:0] _T__7_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_87;
  reg [15:0] _T__7_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_88;
  wire [15:0] _T__7_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_89;
  wire [15:0] _T__7_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__7_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__7_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__7_1__T_17_en_pipe_0;
  reg [31:0] _RAND_90;
  reg [1:0] _T__7_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_91;
  reg [15:0] _T__7_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_92;
  wire [15:0] _T__7_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_93;
  wire [15:0] _T__7_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__7_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__7_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__7_2__T_17_en_pipe_0;
  reg [31:0] _RAND_94;
  reg [1:0] _T__7_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_95;
  reg [15:0] _T__8_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_96;
  wire [15:0] _T__8_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_97;
  wire [15:0] _T__8_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__8_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__8_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__8_0__T_17_en_pipe_0;
  reg [31:0] _RAND_98;
  reg [1:0] _T__8_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_99;
  reg [15:0] _T__8_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_100;
  wire [15:0] _T__8_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_101;
  wire [15:0] _T__8_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__8_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__8_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__8_1__T_17_en_pipe_0;
  reg [31:0] _RAND_102;
  reg [1:0] _T__8_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_103;
  reg [15:0] _T__8_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_104;
  wire [15:0] _T__8_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_105;
  wire [15:0] _T__8_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__8_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__8_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__8_2__T_17_en_pipe_0;
  reg [31:0] _RAND_106;
  reg [1:0] _T__8_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_107;
  reg [15:0] _T__9_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_108;
  wire [15:0] _T__9_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_109;
  wire [15:0] _T__9_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__9_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__9_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__9_0__T_17_en_pipe_0;
  reg [31:0] _RAND_110;
  reg [1:0] _T__9_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_111;
  reg [15:0] _T__9_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_112;
  wire [15:0] _T__9_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_113;
  wire [15:0] _T__9_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__9_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__9_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__9_1__T_17_en_pipe_0;
  reg [31:0] _RAND_114;
  reg [1:0] _T__9_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_115;
  reg [15:0] _T__9_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_116;
  wire [15:0] _T__9_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_117;
  wire [15:0] _T__9_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__9_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__9_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__9_2__T_17_en_pipe_0;
  reg [31:0] _RAND_118;
  reg [1:0] _T__9_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_119;
  reg [15:0] _T__10_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_120;
  wire [15:0] _T__10_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_121;
  wire [15:0] _T__10_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__10_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__10_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__10_0__T_17_en_pipe_0;
  reg [31:0] _RAND_122;
  reg [1:0] _T__10_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_123;
  reg [15:0] _T__10_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_124;
  wire [15:0] _T__10_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_125;
  wire [15:0] _T__10_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__10_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__10_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__10_1__T_17_en_pipe_0;
  reg [31:0] _RAND_126;
  reg [1:0] _T__10_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_127;
  reg [15:0] _T__10_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_128;
  wire [15:0] _T__10_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_129;
  wire [15:0] _T__10_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__10_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__10_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__10_2__T_17_en_pipe_0;
  reg [31:0] _RAND_130;
  reg [1:0] _T__10_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_131;
  reg [15:0] _T__11_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_132;
  wire [15:0] _T__11_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_133;
  wire [15:0] _T__11_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__11_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__11_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__11_0__T_17_en_pipe_0;
  reg [31:0] _RAND_134;
  reg [1:0] _T__11_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_135;
  reg [15:0] _T__11_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_136;
  wire [15:0] _T__11_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_137;
  wire [15:0] _T__11_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__11_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__11_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__11_1__T_17_en_pipe_0;
  reg [31:0] _RAND_138;
  reg [1:0] _T__11_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_139;
  reg [15:0] _T__11_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_140;
  wire [15:0] _T__11_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_141;
  wire [15:0] _T__11_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__11_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__11_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__11_2__T_17_en_pipe_0;
  reg [31:0] _RAND_142;
  reg [1:0] _T__11_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_143;
  reg [15:0] _T__12_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_144;
  wire [15:0] _T__12_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_145;
  wire [15:0] _T__12_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__12_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__12_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__12_0__T_17_en_pipe_0;
  reg [31:0] _RAND_146;
  reg [1:0] _T__12_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_147;
  reg [15:0] _T__12_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_148;
  wire [15:0] _T__12_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_149;
  wire [15:0] _T__12_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__12_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__12_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__12_1__T_17_en_pipe_0;
  reg [31:0] _RAND_150;
  reg [1:0] _T__12_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_151;
  reg [15:0] _T__12_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_152;
  wire [15:0] _T__12_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_153;
  wire [15:0] _T__12_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__12_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__12_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__12_2__T_17_en_pipe_0;
  reg [31:0] _RAND_154;
  reg [1:0] _T__12_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_155;
  reg [15:0] _T__13_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_156;
  wire [15:0] _T__13_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_157;
  wire [15:0] _T__13_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__13_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__13_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__13_0__T_17_en_pipe_0;
  reg [31:0] _RAND_158;
  reg [1:0] _T__13_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_159;
  reg [15:0] _T__13_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_160;
  wire [15:0] _T__13_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_161;
  wire [15:0] _T__13_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__13_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__13_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__13_1__T_17_en_pipe_0;
  reg [31:0] _RAND_162;
  reg [1:0] _T__13_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_163;
  reg [15:0] _T__13_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_164;
  wire [15:0] _T__13_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_165;
  wire [15:0] _T__13_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__13_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__13_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__13_2__T_17_en_pipe_0;
  reg [31:0] _RAND_166;
  reg [1:0] _T__13_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_167;
  reg [15:0] _T__14_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_168;
  wire [15:0] _T__14_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_169;
  wire [15:0] _T__14_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__14_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__14_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__14_0__T_17_en_pipe_0;
  reg [31:0] _RAND_170;
  reg [1:0] _T__14_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_171;
  reg [15:0] _T__14_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_172;
  wire [15:0] _T__14_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_173;
  wire [15:0] _T__14_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__14_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__14_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__14_1__T_17_en_pipe_0;
  reg [31:0] _RAND_174;
  reg [1:0] _T__14_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_175;
  reg [15:0] _T__14_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_176;
  wire [15:0] _T__14_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_177;
  wire [15:0] _T__14_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__14_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__14_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__14_2__T_17_en_pipe_0;
  reg [31:0] _RAND_178;
  reg [1:0] _T__14_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_179;
  reg [15:0] _T__15_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_180;
  wire [15:0] _T__15_0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_181;
  wire [15:0] _T__15_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__15_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__15_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__15_0__T_17_en_pipe_0;
  reg [31:0] _RAND_182;
  reg [1:0] _T__15_0__T_17_addr_pipe_0;
  reg [31:0] _RAND_183;
  reg [15:0] _T__15_1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_184;
  wire [15:0] _T__15_1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_185;
  wire [15:0] _T__15_1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__15_1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__15_1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__15_1__T_17_en_pipe_0;
  reg [31:0] _RAND_186;
  reg [1:0] _T__15_1__T_17_addr_pipe_0;
  reg [31:0] _RAND_187;
  reg [15:0] _T__15_2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_188;
  wire [15:0] _T__15_2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_189;
  wire [15:0] _T__15_2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15_2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__15_2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__15_2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__15_2__T_17_en_pipe_0;
  reg [31:0] _RAND_190;
  reg [1:0] _T__15_2__T_17_addr_pipe_0;
  reg [31:0] _RAND_191;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_192;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_193;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_194;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_11; // @[Counter.scala 38:22]
  wire  _T_12; // @[FIFO.scala 42:39]
  wire  _T_18; // @[Counter.scala 37:24]
  wire [1:0] _T_20; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  wire  _GEN_166; // @[FIFO.scala 39:15]
  assign _T__0_0__T_17_addr = _T__0_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_0__T_17_data = _T__0_0[_T__0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__0_0__T_17_data = _T__0_0__T_17_addr >= 2'h3 ? _RAND_1[15:0] : _T__0_0[_T__0_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_0__T_5_data = I_0_0;
  assign _T__0_0__T_5_addr = value_2;
  assign _T__0_0__T_5_mask = 1'h1;
  assign _T__0_0__T_5_en = valid_up;
  assign _T__0_1__T_17_addr = _T__0_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_1__T_17_data = _T__0_1[_T__0_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__0_1__T_17_data = _T__0_1__T_17_addr >= 2'h3 ? _RAND_5[15:0] : _T__0_1[_T__0_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_1__T_5_data = I_0_1;
  assign _T__0_1__T_5_addr = value_2;
  assign _T__0_1__T_5_mask = 1'h1;
  assign _T__0_1__T_5_en = valid_up;
  assign _T__0_2__T_17_addr = _T__0_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_2__T_17_data = _T__0_2[_T__0_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__0_2__T_17_data = _T__0_2__T_17_addr >= 2'h3 ? _RAND_9[15:0] : _T__0_2[_T__0_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0_2__T_5_data = I_0_2;
  assign _T__0_2__T_5_addr = value_2;
  assign _T__0_2__T_5_mask = 1'h1;
  assign _T__0_2__T_5_en = valid_up;
  assign _T__1_0__T_17_addr = _T__1_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_0__T_17_data = _T__1_0[_T__1_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__1_0__T_17_data = _T__1_0__T_17_addr >= 2'h3 ? _RAND_13[15:0] : _T__1_0[_T__1_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_0__T_5_data = I_1_0;
  assign _T__1_0__T_5_addr = value_2;
  assign _T__1_0__T_5_mask = 1'h1;
  assign _T__1_0__T_5_en = valid_up;
  assign _T__1_1__T_17_addr = _T__1_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_1__T_17_data = _T__1_1[_T__1_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__1_1__T_17_data = _T__1_1__T_17_addr >= 2'h3 ? _RAND_17[15:0] : _T__1_1[_T__1_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_1__T_5_data = I_1_1;
  assign _T__1_1__T_5_addr = value_2;
  assign _T__1_1__T_5_mask = 1'h1;
  assign _T__1_1__T_5_en = valid_up;
  assign _T__1_2__T_17_addr = _T__1_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_2__T_17_data = _T__1_2[_T__1_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__1_2__T_17_data = _T__1_2__T_17_addr >= 2'h3 ? _RAND_21[15:0] : _T__1_2[_T__1_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1_2__T_5_data = I_1_2;
  assign _T__1_2__T_5_addr = value_2;
  assign _T__1_2__T_5_mask = 1'h1;
  assign _T__1_2__T_5_en = valid_up;
  assign _T__2_0__T_17_addr = _T__2_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_0__T_17_data = _T__2_0[_T__2_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__2_0__T_17_data = _T__2_0__T_17_addr >= 2'h3 ? _RAND_25[15:0] : _T__2_0[_T__2_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_0__T_5_data = I_2_0;
  assign _T__2_0__T_5_addr = value_2;
  assign _T__2_0__T_5_mask = 1'h1;
  assign _T__2_0__T_5_en = valid_up;
  assign _T__2_1__T_17_addr = _T__2_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_1__T_17_data = _T__2_1[_T__2_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__2_1__T_17_data = _T__2_1__T_17_addr >= 2'h3 ? _RAND_29[15:0] : _T__2_1[_T__2_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_1__T_5_data = I_2_1;
  assign _T__2_1__T_5_addr = value_2;
  assign _T__2_1__T_5_mask = 1'h1;
  assign _T__2_1__T_5_en = valid_up;
  assign _T__2_2__T_17_addr = _T__2_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_2__T_17_data = _T__2_2[_T__2_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__2_2__T_17_data = _T__2_2__T_17_addr >= 2'h3 ? _RAND_33[15:0] : _T__2_2[_T__2_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2_2__T_5_data = I_2_2;
  assign _T__2_2__T_5_addr = value_2;
  assign _T__2_2__T_5_mask = 1'h1;
  assign _T__2_2__T_5_en = valid_up;
  assign _T__3_0__T_17_addr = _T__3_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_0__T_17_data = _T__3_0[_T__3_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__3_0__T_17_data = _T__3_0__T_17_addr >= 2'h3 ? _RAND_37[15:0] : _T__3_0[_T__3_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_0__T_5_data = I_3_0;
  assign _T__3_0__T_5_addr = value_2;
  assign _T__3_0__T_5_mask = 1'h1;
  assign _T__3_0__T_5_en = valid_up;
  assign _T__3_1__T_17_addr = _T__3_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_1__T_17_data = _T__3_1[_T__3_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__3_1__T_17_data = _T__3_1__T_17_addr >= 2'h3 ? _RAND_41[15:0] : _T__3_1[_T__3_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_1__T_5_data = I_3_1;
  assign _T__3_1__T_5_addr = value_2;
  assign _T__3_1__T_5_mask = 1'h1;
  assign _T__3_1__T_5_en = valid_up;
  assign _T__3_2__T_17_addr = _T__3_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_2__T_17_data = _T__3_2[_T__3_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__3_2__T_17_data = _T__3_2__T_17_addr >= 2'h3 ? _RAND_45[15:0] : _T__3_2[_T__3_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3_2__T_5_data = I_3_2;
  assign _T__3_2__T_5_addr = value_2;
  assign _T__3_2__T_5_mask = 1'h1;
  assign _T__3_2__T_5_en = valid_up;
  assign _T__4_0__T_17_addr = _T__4_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_0__T_17_data = _T__4_0[_T__4_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__4_0__T_17_data = _T__4_0__T_17_addr >= 2'h3 ? _RAND_49[15:0] : _T__4_0[_T__4_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_0__T_5_data = I_4_0;
  assign _T__4_0__T_5_addr = value_2;
  assign _T__4_0__T_5_mask = 1'h1;
  assign _T__4_0__T_5_en = valid_up;
  assign _T__4_1__T_17_addr = _T__4_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_1__T_17_data = _T__4_1[_T__4_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__4_1__T_17_data = _T__4_1__T_17_addr >= 2'h3 ? _RAND_53[15:0] : _T__4_1[_T__4_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_1__T_5_data = I_4_1;
  assign _T__4_1__T_5_addr = value_2;
  assign _T__4_1__T_5_mask = 1'h1;
  assign _T__4_1__T_5_en = valid_up;
  assign _T__4_2__T_17_addr = _T__4_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_2__T_17_data = _T__4_2[_T__4_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__4_2__T_17_data = _T__4_2__T_17_addr >= 2'h3 ? _RAND_57[15:0] : _T__4_2[_T__4_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4_2__T_5_data = I_4_2;
  assign _T__4_2__T_5_addr = value_2;
  assign _T__4_2__T_5_mask = 1'h1;
  assign _T__4_2__T_5_en = valid_up;
  assign _T__5_0__T_17_addr = _T__5_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_0__T_17_data = _T__5_0[_T__5_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__5_0__T_17_data = _T__5_0__T_17_addr >= 2'h3 ? _RAND_61[15:0] : _T__5_0[_T__5_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_0__T_5_data = I_5_0;
  assign _T__5_0__T_5_addr = value_2;
  assign _T__5_0__T_5_mask = 1'h1;
  assign _T__5_0__T_5_en = valid_up;
  assign _T__5_1__T_17_addr = _T__5_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_1__T_17_data = _T__5_1[_T__5_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__5_1__T_17_data = _T__5_1__T_17_addr >= 2'h3 ? _RAND_65[15:0] : _T__5_1[_T__5_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_1__T_5_data = I_5_1;
  assign _T__5_1__T_5_addr = value_2;
  assign _T__5_1__T_5_mask = 1'h1;
  assign _T__5_1__T_5_en = valid_up;
  assign _T__5_2__T_17_addr = _T__5_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_2__T_17_data = _T__5_2[_T__5_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__5_2__T_17_data = _T__5_2__T_17_addr >= 2'h3 ? _RAND_69[15:0] : _T__5_2[_T__5_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5_2__T_5_data = I_5_2;
  assign _T__5_2__T_5_addr = value_2;
  assign _T__5_2__T_5_mask = 1'h1;
  assign _T__5_2__T_5_en = valid_up;
  assign _T__6_0__T_17_addr = _T__6_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_0__T_17_data = _T__6_0[_T__6_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__6_0__T_17_data = _T__6_0__T_17_addr >= 2'h3 ? _RAND_73[15:0] : _T__6_0[_T__6_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_0__T_5_data = I_6_0;
  assign _T__6_0__T_5_addr = value_2;
  assign _T__6_0__T_5_mask = 1'h1;
  assign _T__6_0__T_5_en = valid_up;
  assign _T__6_1__T_17_addr = _T__6_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_1__T_17_data = _T__6_1[_T__6_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__6_1__T_17_data = _T__6_1__T_17_addr >= 2'h3 ? _RAND_77[15:0] : _T__6_1[_T__6_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_1__T_5_data = I_6_1;
  assign _T__6_1__T_5_addr = value_2;
  assign _T__6_1__T_5_mask = 1'h1;
  assign _T__6_1__T_5_en = valid_up;
  assign _T__6_2__T_17_addr = _T__6_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_2__T_17_data = _T__6_2[_T__6_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__6_2__T_17_data = _T__6_2__T_17_addr >= 2'h3 ? _RAND_81[15:0] : _T__6_2[_T__6_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6_2__T_5_data = I_6_2;
  assign _T__6_2__T_5_addr = value_2;
  assign _T__6_2__T_5_mask = 1'h1;
  assign _T__6_2__T_5_en = valid_up;
  assign _T__7_0__T_17_addr = _T__7_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_0__T_17_data = _T__7_0[_T__7_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__7_0__T_17_data = _T__7_0__T_17_addr >= 2'h3 ? _RAND_85[15:0] : _T__7_0[_T__7_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_0__T_5_data = I_7_0;
  assign _T__7_0__T_5_addr = value_2;
  assign _T__7_0__T_5_mask = 1'h1;
  assign _T__7_0__T_5_en = valid_up;
  assign _T__7_1__T_17_addr = _T__7_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_1__T_17_data = _T__7_1[_T__7_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__7_1__T_17_data = _T__7_1__T_17_addr >= 2'h3 ? _RAND_89[15:0] : _T__7_1[_T__7_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_1__T_5_data = I_7_1;
  assign _T__7_1__T_5_addr = value_2;
  assign _T__7_1__T_5_mask = 1'h1;
  assign _T__7_1__T_5_en = valid_up;
  assign _T__7_2__T_17_addr = _T__7_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_2__T_17_data = _T__7_2[_T__7_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__7_2__T_17_data = _T__7_2__T_17_addr >= 2'h3 ? _RAND_93[15:0] : _T__7_2[_T__7_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7_2__T_5_data = I_7_2;
  assign _T__7_2__T_5_addr = value_2;
  assign _T__7_2__T_5_mask = 1'h1;
  assign _T__7_2__T_5_en = valid_up;
  assign _T__8_0__T_17_addr = _T__8_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_0__T_17_data = _T__8_0[_T__8_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__8_0__T_17_data = _T__8_0__T_17_addr >= 2'h3 ? _RAND_97[15:0] : _T__8_0[_T__8_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_0__T_5_data = I_8_0;
  assign _T__8_0__T_5_addr = value_2;
  assign _T__8_0__T_5_mask = 1'h1;
  assign _T__8_0__T_5_en = valid_up;
  assign _T__8_1__T_17_addr = _T__8_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_1__T_17_data = _T__8_1[_T__8_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__8_1__T_17_data = _T__8_1__T_17_addr >= 2'h3 ? _RAND_101[15:0] : _T__8_1[_T__8_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_1__T_5_data = I_8_1;
  assign _T__8_1__T_5_addr = value_2;
  assign _T__8_1__T_5_mask = 1'h1;
  assign _T__8_1__T_5_en = valid_up;
  assign _T__8_2__T_17_addr = _T__8_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_2__T_17_data = _T__8_2[_T__8_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__8_2__T_17_data = _T__8_2__T_17_addr >= 2'h3 ? _RAND_105[15:0] : _T__8_2[_T__8_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8_2__T_5_data = I_8_2;
  assign _T__8_2__T_5_addr = value_2;
  assign _T__8_2__T_5_mask = 1'h1;
  assign _T__8_2__T_5_en = valid_up;
  assign _T__9_0__T_17_addr = _T__9_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_0__T_17_data = _T__9_0[_T__9_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__9_0__T_17_data = _T__9_0__T_17_addr >= 2'h3 ? _RAND_109[15:0] : _T__9_0[_T__9_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_0__T_5_data = I_9_0;
  assign _T__9_0__T_5_addr = value_2;
  assign _T__9_0__T_5_mask = 1'h1;
  assign _T__9_0__T_5_en = valid_up;
  assign _T__9_1__T_17_addr = _T__9_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_1__T_17_data = _T__9_1[_T__9_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__9_1__T_17_data = _T__9_1__T_17_addr >= 2'h3 ? _RAND_113[15:0] : _T__9_1[_T__9_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_1__T_5_data = I_9_1;
  assign _T__9_1__T_5_addr = value_2;
  assign _T__9_1__T_5_mask = 1'h1;
  assign _T__9_1__T_5_en = valid_up;
  assign _T__9_2__T_17_addr = _T__9_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_2__T_17_data = _T__9_2[_T__9_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__9_2__T_17_data = _T__9_2__T_17_addr >= 2'h3 ? _RAND_117[15:0] : _T__9_2[_T__9_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9_2__T_5_data = I_9_2;
  assign _T__9_2__T_5_addr = value_2;
  assign _T__9_2__T_5_mask = 1'h1;
  assign _T__9_2__T_5_en = valid_up;
  assign _T__10_0__T_17_addr = _T__10_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_0__T_17_data = _T__10_0[_T__10_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__10_0__T_17_data = _T__10_0__T_17_addr >= 2'h3 ? _RAND_121[15:0] : _T__10_0[_T__10_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_0__T_5_data = I_10_0;
  assign _T__10_0__T_5_addr = value_2;
  assign _T__10_0__T_5_mask = 1'h1;
  assign _T__10_0__T_5_en = valid_up;
  assign _T__10_1__T_17_addr = _T__10_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_1__T_17_data = _T__10_1[_T__10_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__10_1__T_17_data = _T__10_1__T_17_addr >= 2'h3 ? _RAND_125[15:0] : _T__10_1[_T__10_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_1__T_5_data = I_10_1;
  assign _T__10_1__T_5_addr = value_2;
  assign _T__10_1__T_5_mask = 1'h1;
  assign _T__10_1__T_5_en = valid_up;
  assign _T__10_2__T_17_addr = _T__10_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_2__T_17_data = _T__10_2[_T__10_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__10_2__T_17_data = _T__10_2__T_17_addr >= 2'h3 ? _RAND_129[15:0] : _T__10_2[_T__10_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10_2__T_5_data = I_10_2;
  assign _T__10_2__T_5_addr = value_2;
  assign _T__10_2__T_5_mask = 1'h1;
  assign _T__10_2__T_5_en = valid_up;
  assign _T__11_0__T_17_addr = _T__11_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_0__T_17_data = _T__11_0[_T__11_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__11_0__T_17_data = _T__11_0__T_17_addr >= 2'h3 ? _RAND_133[15:0] : _T__11_0[_T__11_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_0__T_5_data = I_11_0;
  assign _T__11_0__T_5_addr = value_2;
  assign _T__11_0__T_5_mask = 1'h1;
  assign _T__11_0__T_5_en = valid_up;
  assign _T__11_1__T_17_addr = _T__11_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_1__T_17_data = _T__11_1[_T__11_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__11_1__T_17_data = _T__11_1__T_17_addr >= 2'h3 ? _RAND_137[15:0] : _T__11_1[_T__11_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_1__T_5_data = I_11_1;
  assign _T__11_1__T_5_addr = value_2;
  assign _T__11_1__T_5_mask = 1'h1;
  assign _T__11_1__T_5_en = valid_up;
  assign _T__11_2__T_17_addr = _T__11_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_2__T_17_data = _T__11_2[_T__11_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__11_2__T_17_data = _T__11_2__T_17_addr >= 2'h3 ? _RAND_141[15:0] : _T__11_2[_T__11_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11_2__T_5_data = I_11_2;
  assign _T__11_2__T_5_addr = value_2;
  assign _T__11_2__T_5_mask = 1'h1;
  assign _T__11_2__T_5_en = valid_up;
  assign _T__12_0__T_17_addr = _T__12_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_0__T_17_data = _T__12_0[_T__12_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__12_0__T_17_data = _T__12_0__T_17_addr >= 2'h3 ? _RAND_145[15:0] : _T__12_0[_T__12_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_0__T_5_data = I_12_0;
  assign _T__12_0__T_5_addr = value_2;
  assign _T__12_0__T_5_mask = 1'h1;
  assign _T__12_0__T_5_en = valid_up;
  assign _T__12_1__T_17_addr = _T__12_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_1__T_17_data = _T__12_1[_T__12_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__12_1__T_17_data = _T__12_1__T_17_addr >= 2'h3 ? _RAND_149[15:0] : _T__12_1[_T__12_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_1__T_5_data = I_12_1;
  assign _T__12_1__T_5_addr = value_2;
  assign _T__12_1__T_5_mask = 1'h1;
  assign _T__12_1__T_5_en = valid_up;
  assign _T__12_2__T_17_addr = _T__12_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_2__T_17_data = _T__12_2[_T__12_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__12_2__T_17_data = _T__12_2__T_17_addr >= 2'h3 ? _RAND_153[15:0] : _T__12_2[_T__12_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12_2__T_5_data = I_12_2;
  assign _T__12_2__T_5_addr = value_2;
  assign _T__12_2__T_5_mask = 1'h1;
  assign _T__12_2__T_5_en = valid_up;
  assign _T__13_0__T_17_addr = _T__13_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_0__T_17_data = _T__13_0[_T__13_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__13_0__T_17_data = _T__13_0__T_17_addr >= 2'h3 ? _RAND_157[15:0] : _T__13_0[_T__13_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_0__T_5_data = I_13_0;
  assign _T__13_0__T_5_addr = value_2;
  assign _T__13_0__T_5_mask = 1'h1;
  assign _T__13_0__T_5_en = valid_up;
  assign _T__13_1__T_17_addr = _T__13_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_1__T_17_data = _T__13_1[_T__13_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__13_1__T_17_data = _T__13_1__T_17_addr >= 2'h3 ? _RAND_161[15:0] : _T__13_1[_T__13_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_1__T_5_data = I_13_1;
  assign _T__13_1__T_5_addr = value_2;
  assign _T__13_1__T_5_mask = 1'h1;
  assign _T__13_1__T_5_en = valid_up;
  assign _T__13_2__T_17_addr = _T__13_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_2__T_17_data = _T__13_2[_T__13_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__13_2__T_17_data = _T__13_2__T_17_addr >= 2'h3 ? _RAND_165[15:0] : _T__13_2[_T__13_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13_2__T_5_data = I_13_2;
  assign _T__13_2__T_5_addr = value_2;
  assign _T__13_2__T_5_mask = 1'h1;
  assign _T__13_2__T_5_en = valid_up;
  assign _T__14_0__T_17_addr = _T__14_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_0__T_17_data = _T__14_0[_T__14_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__14_0__T_17_data = _T__14_0__T_17_addr >= 2'h3 ? _RAND_169[15:0] : _T__14_0[_T__14_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_0__T_5_data = I_14_0;
  assign _T__14_0__T_5_addr = value_2;
  assign _T__14_0__T_5_mask = 1'h1;
  assign _T__14_0__T_5_en = valid_up;
  assign _T__14_1__T_17_addr = _T__14_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_1__T_17_data = _T__14_1[_T__14_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__14_1__T_17_data = _T__14_1__T_17_addr >= 2'h3 ? _RAND_173[15:0] : _T__14_1[_T__14_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_1__T_5_data = I_14_1;
  assign _T__14_1__T_5_addr = value_2;
  assign _T__14_1__T_5_mask = 1'h1;
  assign _T__14_1__T_5_en = valid_up;
  assign _T__14_2__T_17_addr = _T__14_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_2__T_17_data = _T__14_2[_T__14_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__14_2__T_17_data = _T__14_2__T_17_addr >= 2'h3 ? _RAND_177[15:0] : _T__14_2[_T__14_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14_2__T_5_data = I_14_2;
  assign _T__14_2__T_5_addr = value_2;
  assign _T__14_2__T_5_mask = 1'h1;
  assign _T__14_2__T_5_en = valid_up;
  assign _T__15_0__T_17_addr = _T__15_0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_0__T_17_data = _T__15_0[_T__15_0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__15_0__T_17_data = _T__15_0__T_17_addr >= 2'h3 ? _RAND_181[15:0] : _T__15_0[_T__15_0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_0__T_5_data = I_15_0;
  assign _T__15_0__T_5_addr = value_2;
  assign _T__15_0__T_5_mask = 1'h1;
  assign _T__15_0__T_5_en = valid_up;
  assign _T__15_1__T_17_addr = _T__15_1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_1__T_17_data = _T__15_1[_T__15_1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__15_1__T_17_data = _T__15_1__T_17_addr >= 2'h3 ? _RAND_185[15:0] : _T__15_1[_T__15_1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_1__T_5_data = I_15_1;
  assign _T__15_1__T_5_addr = value_2;
  assign _T__15_1__T_5_mask = 1'h1;
  assign _T__15_1__T_5_en = valid_up;
  assign _T__15_2__T_17_addr = _T__15_2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_2__T_17_data = _T__15_2[_T__15_2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__15_2__T_17_data = _T__15_2__T_17_addr >= 2'h3 ? _RAND_189[15:0] : _T__15_2[_T__15_2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15_2__T_5_data = I_15_2;
  assign _T__15_2__T_5_addr = value_2;
  assign _T__15_2__T_5_mask = 1'h1;
  assign _T__15_2__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_11 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_12 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_18 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_20 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_12 & _T_12; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0 = _T__0_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_0_1 = _T__0_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_0_2 = _T__0_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_1_0 = _T__1_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_1_1 = _T__1_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_1_2 = _T__1_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_2_0 = _T__2_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_2_1 = _T__2_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_2_2 = _T__2_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_3_0 = _T__3_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_3_1 = _T__3_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_3_2 = _T__3_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_4_0 = _T__4_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_4_1 = _T__4_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_4_2 = _T__4_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_5_0 = _T__5_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_5_1 = _T__5_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_5_2 = _T__5_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_6_0 = _T__6_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_6_1 = _T__6_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_6_2 = _T__6_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_7_0 = _T__7_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_7_1 = _T__7_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_7_2 = _T__7_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_8_0 = _T__8_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_8_1 = _T__8_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_8_2 = _T__8_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_9_0 = _T__9_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_9_1 = _T__9_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_9_2 = _T__9_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_10_0 = _T__10_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_10_1 = _T__10_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_10_2 = _T__10_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_11_0 = _T__11_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_11_1 = _T__11_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_11_2 = _T__11_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_12_0 = _T__12_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_12_1 = _T__12_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_12_2 = _T__12_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_13_0 = _T__13_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_13_1 = _T__13_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_13_2 = _T__13_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_14_0 = _T__14_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_14_1 = _T__14_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_14_2 = _T__14_2__T_17_data; // @[FIFO.scala 43:11]
  assign O_15_0 = _T__15_0__T_17_data; // @[FIFO.scala 43:11]
  assign O_15_1 = _T__15_1__T_17_data; // @[FIFO.scala 43:11]
  assign O_15_2 = _T__15_2__T_17_data; // @[FIFO.scala 43:11]
  assign _GEN_166 = valid_up & _T_6; // @[FIFO.scala 39:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__0_0[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0_0__T_17_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__0_0__T_17_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__0_1[initvar] = _RAND_4[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__0_1__T_17_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__0_1__T_17_addr_pipe_0 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__0_2[initvar] = _RAND_8[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__0_2__T_17_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__0_2__T_17_addr_pipe_0 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__1_0[initvar] = _RAND_12[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__1_0__T_17_en_pipe_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__1_0__T_17_addr_pipe_0 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__1_1[initvar] = _RAND_16[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__1_1__T_17_en_pipe_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__1_1__T_17_addr_pipe_0 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__1_2[initvar] = _RAND_20[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__1_2__T_17_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__1_2__T_17_addr_pipe_0 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__2_0[initvar] = _RAND_24[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__2_0__T_17_en_pipe_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__2_0__T_17_addr_pipe_0 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__2_1[initvar] = _RAND_28[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__2_1__T_17_en_pipe_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__2_1__T_17_addr_pipe_0 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__2_2[initvar] = _RAND_32[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__2_2__T_17_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__2_2__T_17_addr_pipe_0 = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__3_0[initvar] = _RAND_36[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_37 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__3_0__T_17_en_pipe_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__3_0__T_17_addr_pipe_0 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__3_1[initvar] = _RAND_40[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_41 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T__3_1__T_17_en_pipe_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T__3_1__T_17_addr_pipe_0 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__3_2[initvar] = _RAND_44[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T__3_2__T_17_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T__3_2__T_17_addr_pipe_0 = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__4_0[initvar] = _RAND_48[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_49 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T__4_0__T_17_en_pipe_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T__4_0__T_17_addr_pipe_0 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__4_1[initvar] = _RAND_52[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_53 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T__4_1__T_17_en_pipe_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T__4_1__T_17_addr_pipe_0 = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__4_2[initvar] = _RAND_56[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T__4_2__T_17_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T__4_2__T_17_addr_pipe_0 = _RAND_59[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__5_0[initvar] = _RAND_60[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_61 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T__5_0__T_17_en_pipe_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T__5_0__T_17_addr_pipe_0 = _RAND_63[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__5_1[initvar] = _RAND_64[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_65 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T__5_1__T_17_en_pipe_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T__5_1__T_17_addr_pipe_0 = _RAND_67[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__5_2[initvar] = _RAND_68[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_69 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T__5_2__T_17_en_pipe_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T__5_2__T_17_addr_pipe_0 = _RAND_71[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__6_0[initvar] = _RAND_72[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_73 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T__6_0__T_17_en_pipe_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T__6_0__T_17_addr_pipe_0 = _RAND_75[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__6_1[initvar] = _RAND_76[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_77 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T__6_1__T_17_en_pipe_0 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T__6_1__T_17_addr_pipe_0 = _RAND_79[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__6_2[initvar] = _RAND_80[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_81 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T__6_2__T_17_en_pipe_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T__6_2__T_17_addr_pipe_0 = _RAND_83[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__7_0[initvar] = _RAND_84[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_85 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T__7_0__T_17_en_pipe_0 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T__7_0__T_17_addr_pipe_0 = _RAND_87[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__7_1[initvar] = _RAND_88[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_89 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T__7_1__T_17_en_pipe_0 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T__7_1__T_17_addr_pipe_0 = _RAND_91[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__7_2[initvar] = _RAND_92[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_93 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T__7_2__T_17_en_pipe_0 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T__7_2__T_17_addr_pipe_0 = _RAND_95[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__8_0[initvar] = _RAND_96[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_97 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T__8_0__T_17_en_pipe_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T__8_0__T_17_addr_pipe_0 = _RAND_99[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__8_1[initvar] = _RAND_100[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_101 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T__8_1__T_17_en_pipe_0 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T__8_1__T_17_addr_pipe_0 = _RAND_103[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__8_2[initvar] = _RAND_104[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_105 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T__8_2__T_17_en_pipe_0 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T__8_2__T_17_addr_pipe_0 = _RAND_107[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__9_0[initvar] = _RAND_108[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_109 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T__9_0__T_17_en_pipe_0 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T__9_0__T_17_addr_pipe_0 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__9_1[initvar] = _RAND_112[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_113 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T__9_1__T_17_en_pipe_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T__9_1__T_17_addr_pipe_0 = _RAND_115[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__9_2[initvar] = _RAND_116[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_117 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T__9_2__T_17_en_pipe_0 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T__9_2__T_17_addr_pipe_0 = _RAND_119[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__10_0[initvar] = _RAND_120[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_121 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T__10_0__T_17_en_pipe_0 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T__10_0__T_17_addr_pipe_0 = _RAND_123[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__10_1[initvar] = _RAND_124[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_125 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T__10_1__T_17_en_pipe_0 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T__10_1__T_17_addr_pipe_0 = _RAND_127[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__10_2[initvar] = _RAND_128[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_129 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T__10_2__T_17_en_pipe_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T__10_2__T_17_addr_pipe_0 = _RAND_131[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__11_0[initvar] = _RAND_132[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_133 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T__11_0__T_17_en_pipe_0 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T__11_0__T_17_addr_pipe_0 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__11_1[initvar] = _RAND_136[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_137 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T__11_1__T_17_en_pipe_0 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T__11_1__T_17_addr_pipe_0 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__11_2[initvar] = _RAND_140[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_141 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T__11_2__T_17_en_pipe_0 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T__11_2__T_17_addr_pipe_0 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__12_0[initvar] = _RAND_144[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_145 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T__12_0__T_17_en_pipe_0 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T__12_0__T_17_addr_pipe_0 = _RAND_147[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__12_1[initvar] = _RAND_148[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_149 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T__12_1__T_17_en_pipe_0 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T__12_1__T_17_addr_pipe_0 = _RAND_151[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__12_2[initvar] = _RAND_152[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_153 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T__12_2__T_17_en_pipe_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T__12_2__T_17_addr_pipe_0 = _RAND_155[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__13_0[initvar] = _RAND_156[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_157 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T__13_0__T_17_en_pipe_0 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T__13_0__T_17_addr_pipe_0 = _RAND_159[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__13_1[initvar] = _RAND_160[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_161 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T__13_1__T_17_en_pipe_0 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T__13_1__T_17_addr_pipe_0 = _RAND_163[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__13_2[initvar] = _RAND_164[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_165 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T__13_2__T_17_en_pipe_0 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T__13_2__T_17_addr_pipe_0 = _RAND_167[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__14_0[initvar] = _RAND_168[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_169 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T__14_0__T_17_en_pipe_0 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T__14_0__T_17_addr_pipe_0 = _RAND_171[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__14_1[initvar] = _RAND_172[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_173 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T__14_1__T_17_en_pipe_0 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T__14_1__T_17_addr_pipe_0 = _RAND_175[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__14_2[initvar] = _RAND_176[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_177 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T__14_2__T_17_en_pipe_0 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T__14_2__T_17_addr_pipe_0 = _RAND_179[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__15_0[initvar] = _RAND_180[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_181 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T__15_0__T_17_en_pipe_0 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T__15_0__T_17_addr_pipe_0 = _RAND_183[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__15_1[initvar] = _RAND_184[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_185 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T__15_1__T_17_en_pipe_0 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T__15_1__T_17_addr_pipe_0 = _RAND_187[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__15_2[initvar] = _RAND_188[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_189 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T__15_2__T_17_en_pipe_0 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T__15_2__T_17_addr_pipe_0 = _RAND_191[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  value = _RAND_192[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  value_1 = _RAND_193[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  value_2 = _RAND_194[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__0_0__T_5_en & _T__0_0__T_5_mask) begin
      _T__0_0[_T__0_0__T_5_addr] <= _T__0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__0_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__0_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__0_1__T_5_en & _T__0_1__T_5_mask) begin
      _T__0_1[_T__0_1__T_5_addr] <= _T__0_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__0_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__0_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__0_2__T_5_en & _T__0_2__T_5_mask) begin
      _T__0_2[_T__0_2__T_5_addr] <= _T__0_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__0_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__0_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__1_0__T_5_en & _T__1_0__T_5_mask) begin
      _T__1_0[_T__1_0__T_5_addr] <= _T__1_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__1_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__1_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__1_1__T_5_en & _T__1_1__T_5_mask) begin
      _T__1_1[_T__1_1__T_5_addr] <= _T__1_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__1_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__1_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__1_2__T_5_en & _T__1_2__T_5_mask) begin
      _T__1_2[_T__1_2__T_5_addr] <= _T__1_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__1_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__1_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__2_0__T_5_en & _T__2_0__T_5_mask) begin
      _T__2_0[_T__2_0__T_5_addr] <= _T__2_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__2_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__2_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__2_1__T_5_en & _T__2_1__T_5_mask) begin
      _T__2_1[_T__2_1__T_5_addr] <= _T__2_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__2_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__2_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__2_2__T_5_en & _T__2_2__T_5_mask) begin
      _T__2_2[_T__2_2__T_5_addr] <= _T__2_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__2_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__2_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__3_0__T_5_en & _T__3_0__T_5_mask) begin
      _T__3_0[_T__3_0__T_5_addr] <= _T__3_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__3_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__3_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__3_1__T_5_en & _T__3_1__T_5_mask) begin
      _T__3_1[_T__3_1__T_5_addr] <= _T__3_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__3_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__3_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__3_2__T_5_en & _T__3_2__T_5_mask) begin
      _T__3_2[_T__3_2__T_5_addr] <= _T__3_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__3_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__3_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__4_0__T_5_en & _T__4_0__T_5_mask) begin
      _T__4_0[_T__4_0__T_5_addr] <= _T__4_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__4_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__4_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__4_1__T_5_en & _T__4_1__T_5_mask) begin
      _T__4_1[_T__4_1__T_5_addr] <= _T__4_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__4_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__4_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__4_2__T_5_en & _T__4_2__T_5_mask) begin
      _T__4_2[_T__4_2__T_5_addr] <= _T__4_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__4_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__4_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__5_0__T_5_en & _T__5_0__T_5_mask) begin
      _T__5_0[_T__5_0__T_5_addr] <= _T__5_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__5_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__5_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__5_1__T_5_en & _T__5_1__T_5_mask) begin
      _T__5_1[_T__5_1__T_5_addr] <= _T__5_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__5_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__5_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__5_2__T_5_en & _T__5_2__T_5_mask) begin
      _T__5_2[_T__5_2__T_5_addr] <= _T__5_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__5_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__5_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__6_0__T_5_en & _T__6_0__T_5_mask) begin
      _T__6_0[_T__6_0__T_5_addr] <= _T__6_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__6_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__6_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__6_1__T_5_en & _T__6_1__T_5_mask) begin
      _T__6_1[_T__6_1__T_5_addr] <= _T__6_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__6_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__6_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__6_2__T_5_en & _T__6_2__T_5_mask) begin
      _T__6_2[_T__6_2__T_5_addr] <= _T__6_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__6_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__6_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__7_0__T_5_en & _T__7_0__T_5_mask) begin
      _T__7_0[_T__7_0__T_5_addr] <= _T__7_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__7_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__7_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__7_1__T_5_en & _T__7_1__T_5_mask) begin
      _T__7_1[_T__7_1__T_5_addr] <= _T__7_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__7_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__7_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__7_2__T_5_en & _T__7_2__T_5_mask) begin
      _T__7_2[_T__7_2__T_5_addr] <= _T__7_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__7_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__7_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__8_0__T_5_en & _T__8_0__T_5_mask) begin
      _T__8_0[_T__8_0__T_5_addr] <= _T__8_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__8_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__8_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__8_1__T_5_en & _T__8_1__T_5_mask) begin
      _T__8_1[_T__8_1__T_5_addr] <= _T__8_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__8_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__8_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__8_2__T_5_en & _T__8_2__T_5_mask) begin
      _T__8_2[_T__8_2__T_5_addr] <= _T__8_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__8_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__8_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__9_0__T_5_en & _T__9_0__T_5_mask) begin
      _T__9_0[_T__9_0__T_5_addr] <= _T__9_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__9_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__9_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__9_1__T_5_en & _T__9_1__T_5_mask) begin
      _T__9_1[_T__9_1__T_5_addr] <= _T__9_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__9_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__9_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__9_2__T_5_en & _T__9_2__T_5_mask) begin
      _T__9_2[_T__9_2__T_5_addr] <= _T__9_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__9_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__9_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__10_0__T_5_en & _T__10_0__T_5_mask) begin
      _T__10_0[_T__10_0__T_5_addr] <= _T__10_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__10_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__10_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__10_1__T_5_en & _T__10_1__T_5_mask) begin
      _T__10_1[_T__10_1__T_5_addr] <= _T__10_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__10_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__10_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__10_2__T_5_en & _T__10_2__T_5_mask) begin
      _T__10_2[_T__10_2__T_5_addr] <= _T__10_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__10_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__10_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__11_0__T_5_en & _T__11_0__T_5_mask) begin
      _T__11_0[_T__11_0__T_5_addr] <= _T__11_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__11_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__11_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__11_1__T_5_en & _T__11_1__T_5_mask) begin
      _T__11_1[_T__11_1__T_5_addr] <= _T__11_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__11_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__11_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__11_2__T_5_en & _T__11_2__T_5_mask) begin
      _T__11_2[_T__11_2__T_5_addr] <= _T__11_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__11_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__11_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__12_0__T_5_en & _T__12_0__T_5_mask) begin
      _T__12_0[_T__12_0__T_5_addr] <= _T__12_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__12_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__12_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__12_1__T_5_en & _T__12_1__T_5_mask) begin
      _T__12_1[_T__12_1__T_5_addr] <= _T__12_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__12_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__12_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__12_2__T_5_en & _T__12_2__T_5_mask) begin
      _T__12_2[_T__12_2__T_5_addr] <= _T__12_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__12_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__12_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__13_0__T_5_en & _T__13_0__T_5_mask) begin
      _T__13_0[_T__13_0__T_5_addr] <= _T__13_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__13_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__13_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__13_1__T_5_en & _T__13_1__T_5_mask) begin
      _T__13_1[_T__13_1__T_5_addr] <= _T__13_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__13_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__13_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__13_2__T_5_en & _T__13_2__T_5_mask) begin
      _T__13_2[_T__13_2__T_5_addr] <= _T__13_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__13_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__13_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__14_0__T_5_en & _T__14_0__T_5_mask) begin
      _T__14_0[_T__14_0__T_5_addr] <= _T__14_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__14_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__14_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__14_1__T_5_en & _T__14_1__T_5_mask) begin
      _T__14_1[_T__14_1__T_5_addr] <= _T__14_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__14_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__14_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__14_2__T_5_en & _T__14_2__T_5_mask) begin
      _T__14_2[_T__14_2__T_5_addr] <= _T__14_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__14_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__14_2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__15_0__T_5_en & _T__15_0__T_5_mask) begin
      _T__15_0[_T__15_0__T_5_addr] <= _T__15_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__15_0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__15_0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__15_1__T_5_en & _T__15_1__T_5_mask) begin
      _T__15_1[_T__15_1__T_5_addr] <= _T__15_1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__15_1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__15_1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__15_2__T_5_en & _T__15_2__T_5_mask) begin
      _T__15_2[_T__15_2__T_5_addr] <= _T__15_2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__15_2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__15_2__T_17_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_11;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_12) begin
        if (_T_18) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_20;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & ~reset) begin
          $fwrite(32'h80000002,"idc inc\n"); // @[FIFO.scala 39:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SSeqTupleAppender_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I1_0,
  input  [15:0] I1_1,
  input  [15:0] I1_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0_0,
  input  [15:0] I0_0_0_1,
  input  [15:0] I0_0_0_2,
  input  [15:0] I0_0_1_0,
  input  [15:0] I0_0_1_1,
  input  [15:0] I0_0_1_2,
  input  [15:0] I0_1_0_0,
  input  [15:0] I0_1_0_1,
  input  [15:0] I0_1_0_2,
  input  [15:0] I0_1_1_0,
  input  [15:0] I0_1_1_1,
  input  [15:0] I0_1_1_2,
  input  [15:0] I0_2_0_0,
  input  [15:0] I0_2_0_1,
  input  [15:0] I0_2_0_2,
  input  [15:0] I0_2_1_0,
  input  [15:0] I0_2_1_1,
  input  [15:0] I0_2_1_2,
  input  [15:0] I0_3_0_0,
  input  [15:0] I0_3_0_1,
  input  [15:0] I0_3_0_2,
  input  [15:0] I0_3_1_0,
  input  [15:0] I0_3_1_1,
  input  [15:0] I0_3_1_2,
  input  [15:0] I0_4_0_0,
  input  [15:0] I0_4_0_1,
  input  [15:0] I0_4_0_2,
  input  [15:0] I0_4_1_0,
  input  [15:0] I0_4_1_1,
  input  [15:0] I0_4_1_2,
  input  [15:0] I0_5_0_0,
  input  [15:0] I0_5_0_1,
  input  [15:0] I0_5_0_2,
  input  [15:0] I0_5_1_0,
  input  [15:0] I0_5_1_1,
  input  [15:0] I0_5_1_2,
  input  [15:0] I0_6_0_0,
  input  [15:0] I0_6_0_1,
  input  [15:0] I0_6_0_2,
  input  [15:0] I0_6_1_0,
  input  [15:0] I0_6_1_1,
  input  [15:0] I0_6_1_2,
  input  [15:0] I0_7_0_0,
  input  [15:0] I0_7_0_1,
  input  [15:0] I0_7_0_2,
  input  [15:0] I0_7_1_0,
  input  [15:0] I0_7_1_1,
  input  [15:0] I0_7_1_2,
  input  [15:0] I0_8_0_0,
  input  [15:0] I0_8_0_1,
  input  [15:0] I0_8_0_2,
  input  [15:0] I0_8_1_0,
  input  [15:0] I0_8_1_1,
  input  [15:0] I0_8_1_2,
  input  [15:0] I0_9_0_0,
  input  [15:0] I0_9_0_1,
  input  [15:0] I0_9_0_2,
  input  [15:0] I0_9_1_0,
  input  [15:0] I0_9_1_1,
  input  [15:0] I0_9_1_2,
  input  [15:0] I0_10_0_0,
  input  [15:0] I0_10_0_1,
  input  [15:0] I0_10_0_2,
  input  [15:0] I0_10_1_0,
  input  [15:0] I0_10_1_1,
  input  [15:0] I0_10_1_2,
  input  [15:0] I0_11_0_0,
  input  [15:0] I0_11_0_1,
  input  [15:0] I0_11_0_2,
  input  [15:0] I0_11_1_0,
  input  [15:0] I0_11_1_1,
  input  [15:0] I0_11_1_2,
  input  [15:0] I0_12_0_0,
  input  [15:0] I0_12_0_1,
  input  [15:0] I0_12_0_2,
  input  [15:0] I0_12_1_0,
  input  [15:0] I0_12_1_1,
  input  [15:0] I0_12_1_2,
  input  [15:0] I0_13_0_0,
  input  [15:0] I0_13_0_1,
  input  [15:0] I0_13_0_2,
  input  [15:0] I0_13_1_0,
  input  [15:0] I0_13_1_1,
  input  [15:0] I0_13_1_2,
  input  [15:0] I0_14_0_0,
  input  [15:0] I0_14_0_1,
  input  [15:0] I0_14_0_2,
  input  [15:0] I0_14_1_0,
  input  [15:0] I0_14_1_1,
  input  [15:0] I0_14_1_2,
  input  [15:0] I0_15_0_0,
  input  [15:0] I0_15_0_1,
  input  [15:0] I0_15_0_2,
  input  [15:0] I0_15_1_0,
  input  [15:0] I0_15_1_1,
  input  [15:0] I0_15_1_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  input  [15:0] I1_8_0,
  input  [15:0] I1_8_1,
  input  [15:0] I1_8_2,
  input  [15:0] I1_9_0,
  input  [15:0] I1_9_1,
  input  [15:0] I1_9_2,
  input  [15:0] I1_10_0,
  input  [15:0] I1_10_1,
  input  [15:0] I1_10_2,
  input  [15:0] I1_11_0,
  input  [15:0] I1_11_1,
  input  [15:0] I1_11_2,
  input  [15:0] I1_12_0,
  input  [15:0] I1_12_1,
  input  [15:0] I1_12_2,
  input  [15:0] I1_13_0,
  input  [15:0] I1_13_1,
  input  [15:0] I1_13_2,
  input  [15:0] I1_14_0,
  input  [15:0] I1_14_1,
  input  [15:0] I1_14_2,
  input  [15:0] I1_15_0,
  input  [15:0] I1_15_1,
  input  [15:0] I1_15_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_8_1_0,
  output [15:0] O_8_1_1,
  output [15:0] O_8_1_2,
  output [15:0] O_8_2_0,
  output [15:0] O_8_2_1,
  output [15:0] O_8_2_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_9_1_0,
  output [15:0] O_9_1_1,
  output [15:0] O_9_1_2,
  output [15:0] O_9_2_0,
  output [15:0] O_9_2_1,
  output [15:0] O_9_2_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_10_1_0,
  output [15:0] O_10_1_1,
  output [15:0] O_10_1_2,
  output [15:0] O_10_2_0,
  output [15:0] O_10_2_1,
  output [15:0] O_10_2_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_11_1_0,
  output [15:0] O_11_1_1,
  output [15:0] O_11_1_2,
  output [15:0] O_11_2_0,
  output [15:0] O_11_2_1,
  output [15:0] O_11_2_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_12_1_0,
  output [15:0] O_12_1_1,
  output [15:0] O_12_1_2,
  output [15:0] O_12_2_0,
  output [15:0] O_12_2_1,
  output [15:0] O_12_2_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_13_1_0,
  output [15:0] O_13_1_1,
  output [15:0] O_13_1_2,
  output [15:0] O_13_2_0,
  output [15:0] O_13_2_1,
  output [15:0] O_13_2_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_14_1_0,
  output [15:0] O_14_1_1,
  output [15:0] O_14_1_2,
  output [15:0] O_14_2_0,
  output [15:0] O_14_2_1,
  output [15:0] O_14_2_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2,
  output [15:0] O_15_1_0,
  output [15:0] O_15_1_1,
  output [15:0] O_15_1_2,
  output [15:0] O_15_2_0,
  output [15:0] O_15_2_1,
  output [15:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_2_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_3_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_4_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_5_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_6_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_7_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_8_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_9_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_10_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_11_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_12_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_13_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I0_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_2_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_2_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_14_O_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I0_0_1(other_ops_7_I0_0_1),
    .I0_0_2(other_ops_7_I0_0_2),
    .I0_1_0(other_ops_7_I0_1_0),
    .I0_1_1(other_ops_7_I0_1_1),
    .I0_1_2(other_ops_7_I0_1_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I0_0_1(other_ops_8_I0_0_1),
    .I0_0_2(other_ops_8_I0_0_2),
    .I0_1_0(other_ops_8_I0_1_0),
    .I0_1_1(other_ops_8_I0_1_1),
    .I0_1_2(other_ops_8_I0_1_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I0_0_1(other_ops_9_I0_0_1),
    .I0_0_2(other_ops_9_I0_0_2),
    .I0_1_0(other_ops_9_I0_1_0),
    .I0_1_1(other_ops_9_I0_1_1),
    .I0_1_2(other_ops_9_I0_1_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I0_0_1(other_ops_10_I0_0_1),
    .I0_0_2(other_ops_10_I0_0_2),
    .I0_1_0(other_ops_10_I0_1_0),
    .I0_1_1(other_ops_10_I0_1_1),
    .I0_1_2(other_ops_10_I0_1_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I0_0_1(other_ops_11_I0_0_1),
    .I0_0_2(other_ops_11_I0_0_2),
    .I0_1_0(other_ops_11_I0_1_0),
    .I0_1_1(other_ops_11_I0_1_1),
    .I0_1_2(other_ops_11_I0_1_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I0_0_1(other_ops_12_I0_0_1),
    .I0_0_2(other_ops_12_I0_0_2),
    .I0_1_0(other_ops_12_I0_1_0),
    .I0_1_1(other_ops_12_I0_1_1),
    .I0_1_2(other_ops_12_I0_1_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I0_0_1(other_ops_13_I0_0_1),
    .I0_0_2(other_ops_13_I0_0_2),
    .I0_1_0(other_ops_13_I0_1_0),
    .I0_1_1(other_ops_13_I0_1_1),
    .I0_1_2(other_ops_13_I0_1_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I0_0_1(other_ops_14_I0_0_1),
    .I0_0_2(other_ops_14_I0_0_2),
    .I0_1_0(other_ops_14_I0_1_0),
    .I0_1_1(other_ops_14_I0_1_1),
    .I0_1_2(other_ops_14_I0_1_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[Map2S.scala 24:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[Map2S.scala 24:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[Map2S.scala 24:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[Map2S.scala 24:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[Map2S.scala 24:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[Map2S.scala 24:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[Map2S.scala 24:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[Map2S.scala 24:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[Map2S.scala 24:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[Map2S.scala 24:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[Map2S.scala 24:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[Map2S.scala 24:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[Map2S.scala 24:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[Map2S.scala 24:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[Map2S.scala 24:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[Map2S.scala 24:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[Map2S.scala 24:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[Map2S.scala 24:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[Map2S.scala 24:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[Map2S.scala 24:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[Map2S.scala 24:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[Map2S.scala 24:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[Map2S.scala 24:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[Map2S.scala 24:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[Map2S.scala 24:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[Map2S.scala 24:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[Map2S.scala 24:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[Map2S.scala 24:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1 = I0_8_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_2 = I0_8_0_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_0 = I0_8_1_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_1 = I0_8_1_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_2 = I0_8_1_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1 = I0_9_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_2 = I0_9_0_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_0 = I0_9_1_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_1 = I0_9_1_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_2 = I0_9_1_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1 = I0_10_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_2 = I0_10_0_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_0 = I0_10_1_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_1 = I0_10_1_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_2 = I0_10_1_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1 = I0_11_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_2 = I0_11_0_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_0 = I0_11_1_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_1 = I0_11_1_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_2 = I0_11_1_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1 = I0_12_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_2 = I0_12_0_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_0 = I0_12_1_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_1 = I0_12_1_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_2 = I0_12_1_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1 = I0_13_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_2 = I0_13_0_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_0 = I0_13_1_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_1 = I0_13_1_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_2 = I0_13_1_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1 = I0_14_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_2 = I0_14_0_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_0 = I0_14_1_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_1 = I0_14_1_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_2 = I0_14_1_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1 = I0_15_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_2 = I0_15_0_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_0 = I0_15_1_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_1 = I0_15_1_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_2 = I0_15_1_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0_0,
  input  [15:0] I0_0_0_1,
  input  [15:0] I0_0_0_2,
  input  [15:0] I0_0_1_0,
  input  [15:0] I0_0_1_1,
  input  [15:0] I0_0_1_2,
  input  [15:0] I0_1_0_0,
  input  [15:0] I0_1_0_1,
  input  [15:0] I0_1_0_2,
  input  [15:0] I0_1_1_0,
  input  [15:0] I0_1_1_1,
  input  [15:0] I0_1_1_2,
  input  [15:0] I0_2_0_0,
  input  [15:0] I0_2_0_1,
  input  [15:0] I0_2_0_2,
  input  [15:0] I0_2_1_0,
  input  [15:0] I0_2_1_1,
  input  [15:0] I0_2_1_2,
  input  [15:0] I0_3_0_0,
  input  [15:0] I0_3_0_1,
  input  [15:0] I0_3_0_2,
  input  [15:0] I0_3_1_0,
  input  [15:0] I0_3_1_1,
  input  [15:0] I0_3_1_2,
  input  [15:0] I0_4_0_0,
  input  [15:0] I0_4_0_1,
  input  [15:0] I0_4_0_2,
  input  [15:0] I0_4_1_0,
  input  [15:0] I0_4_1_1,
  input  [15:0] I0_4_1_2,
  input  [15:0] I0_5_0_0,
  input  [15:0] I0_5_0_1,
  input  [15:0] I0_5_0_2,
  input  [15:0] I0_5_1_0,
  input  [15:0] I0_5_1_1,
  input  [15:0] I0_5_1_2,
  input  [15:0] I0_6_0_0,
  input  [15:0] I0_6_0_1,
  input  [15:0] I0_6_0_2,
  input  [15:0] I0_6_1_0,
  input  [15:0] I0_6_1_1,
  input  [15:0] I0_6_1_2,
  input  [15:0] I0_7_0_0,
  input  [15:0] I0_7_0_1,
  input  [15:0] I0_7_0_2,
  input  [15:0] I0_7_1_0,
  input  [15:0] I0_7_1_1,
  input  [15:0] I0_7_1_2,
  input  [15:0] I0_8_0_0,
  input  [15:0] I0_8_0_1,
  input  [15:0] I0_8_0_2,
  input  [15:0] I0_8_1_0,
  input  [15:0] I0_8_1_1,
  input  [15:0] I0_8_1_2,
  input  [15:0] I0_9_0_0,
  input  [15:0] I0_9_0_1,
  input  [15:0] I0_9_0_2,
  input  [15:0] I0_9_1_0,
  input  [15:0] I0_9_1_1,
  input  [15:0] I0_9_1_2,
  input  [15:0] I0_10_0_0,
  input  [15:0] I0_10_0_1,
  input  [15:0] I0_10_0_2,
  input  [15:0] I0_10_1_0,
  input  [15:0] I0_10_1_1,
  input  [15:0] I0_10_1_2,
  input  [15:0] I0_11_0_0,
  input  [15:0] I0_11_0_1,
  input  [15:0] I0_11_0_2,
  input  [15:0] I0_11_1_0,
  input  [15:0] I0_11_1_1,
  input  [15:0] I0_11_1_2,
  input  [15:0] I0_12_0_0,
  input  [15:0] I0_12_0_1,
  input  [15:0] I0_12_0_2,
  input  [15:0] I0_12_1_0,
  input  [15:0] I0_12_1_1,
  input  [15:0] I0_12_1_2,
  input  [15:0] I0_13_0_0,
  input  [15:0] I0_13_0_1,
  input  [15:0] I0_13_0_2,
  input  [15:0] I0_13_1_0,
  input  [15:0] I0_13_1_1,
  input  [15:0] I0_13_1_2,
  input  [15:0] I0_14_0_0,
  input  [15:0] I0_14_0_1,
  input  [15:0] I0_14_0_2,
  input  [15:0] I0_14_1_0,
  input  [15:0] I0_14_1_1,
  input  [15:0] I0_14_1_2,
  input  [15:0] I0_15_0_0,
  input  [15:0] I0_15_0_1,
  input  [15:0] I0_15_0_2,
  input  [15:0] I0_15_1_0,
  input  [15:0] I0_15_1_1,
  input  [15:0] I0_15_1_2,
  input  [15:0] I1_0_0,
  input  [15:0] I1_0_1,
  input  [15:0] I1_0_2,
  input  [15:0] I1_1_0,
  input  [15:0] I1_1_1,
  input  [15:0] I1_1_2,
  input  [15:0] I1_2_0,
  input  [15:0] I1_2_1,
  input  [15:0] I1_2_2,
  input  [15:0] I1_3_0,
  input  [15:0] I1_3_1,
  input  [15:0] I1_3_2,
  input  [15:0] I1_4_0,
  input  [15:0] I1_4_1,
  input  [15:0] I1_4_2,
  input  [15:0] I1_5_0,
  input  [15:0] I1_5_1,
  input  [15:0] I1_5_2,
  input  [15:0] I1_6_0,
  input  [15:0] I1_6_1,
  input  [15:0] I1_6_2,
  input  [15:0] I1_7_0,
  input  [15:0] I1_7_1,
  input  [15:0] I1_7_2,
  input  [15:0] I1_8_0,
  input  [15:0] I1_8_1,
  input  [15:0] I1_8_2,
  input  [15:0] I1_9_0,
  input  [15:0] I1_9_1,
  input  [15:0] I1_9_2,
  input  [15:0] I1_10_0,
  input  [15:0] I1_10_1,
  input  [15:0] I1_10_2,
  input  [15:0] I1_11_0,
  input  [15:0] I1_11_1,
  input  [15:0] I1_11_2,
  input  [15:0] I1_12_0,
  input  [15:0] I1_12_1,
  input  [15:0] I1_12_2,
  input  [15:0] I1_13_0,
  input  [15:0] I1_13_1,
  input  [15:0] I1_13_2,
  input  [15:0] I1_14_0,
  input  [15:0] I1_14_1,
  input  [15:0] I1_14_2,
  input  [15:0] I1_15_0,
  input  [15:0] I1_15_1,
  input  [15:0] I1_15_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_8_1_0,
  output [15:0] O_8_1_1,
  output [15:0] O_8_1_2,
  output [15:0] O_8_2_0,
  output [15:0] O_8_2_1,
  output [15:0] O_8_2_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_9_1_0,
  output [15:0] O_9_1_1,
  output [15:0] O_9_1_2,
  output [15:0] O_9_2_0,
  output [15:0] O_9_2_1,
  output [15:0] O_9_2_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_10_1_0,
  output [15:0] O_10_1_1,
  output [15:0] O_10_1_2,
  output [15:0] O_10_2_0,
  output [15:0] O_10_2_1,
  output [15:0] O_10_2_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_11_1_0,
  output [15:0] O_11_1_1,
  output [15:0] O_11_1_2,
  output [15:0] O_11_2_0,
  output [15:0] O_11_2_1,
  output [15:0] O_11_2_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_12_1_0,
  output [15:0] O_12_1_1,
  output [15:0] O_12_1_2,
  output [15:0] O_12_2_0,
  output [15:0] O_12_2_1,
  output [15:0] O_12_2_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_13_1_0,
  output [15:0] O_13_1_1,
  output [15:0] O_13_1_2,
  output [15:0] O_13_2_0,
  output [15:0] O_13_2_1,
  output [15:0] O_13_2_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_14_1_0,
  output [15:0] O_14_1_1,
  output [15:0] O_14_1_2,
  output [15:0] O_14_2_0,
  output [15:0] O_14_2_1,
  output [15:0] O_14_2_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2,
  output [15:0] O_15_1_0,
  output [15:0] O_15_1_1,
  output [15:0] O_15_1_2,
  output [15:0] O_15_2_0,
  output [15:0] O_15_2_1,
  output [15:0] O_15_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_4_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_5_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_6_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_7_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_8_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_9_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_10_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_11_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_12_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_13_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_14_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I0_15_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_8_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_9_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_10_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_11_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_12_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_13_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_14_2; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15_0; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15_1; // @[Map2T.scala 8:20]
  wire [15:0] op_I1_15_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_0_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_1_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_2_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_3_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_4_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_5_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_6_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_7_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_8_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_9_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_10_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_11_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_12_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_13_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_14_2_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_0_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_1_2; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_2_0; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_2_1; // @[Map2T.scala 8:20]
  wire [15:0] op_O_15_2_2; // @[Map2T.scala 8:20]
  Map2S_7 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_4_1_0(op_I0_4_1_0),
    .I0_4_1_1(op_I0_4_1_1),
    .I0_4_1_2(op_I0_4_1_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_5_1_0(op_I0_5_1_0),
    .I0_5_1_1(op_I0_5_1_1),
    .I0_5_1_2(op_I0_5_1_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_6_1_0(op_I0_6_1_0),
    .I0_6_1_1(op_I0_6_1_1),
    .I0_6_1_2(op_I0_6_1_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_7_1_0(op_I0_7_1_0),
    .I0_7_1_1(op_I0_7_1_1),
    .I0_7_1_2(op_I0_7_1_2),
    .I0_8_0_0(op_I0_8_0_0),
    .I0_8_0_1(op_I0_8_0_1),
    .I0_8_0_2(op_I0_8_0_2),
    .I0_8_1_0(op_I0_8_1_0),
    .I0_8_1_1(op_I0_8_1_1),
    .I0_8_1_2(op_I0_8_1_2),
    .I0_9_0_0(op_I0_9_0_0),
    .I0_9_0_1(op_I0_9_0_1),
    .I0_9_0_2(op_I0_9_0_2),
    .I0_9_1_0(op_I0_9_1_0),
    .I0_9_1_1(op_I0_9_1_1),
    .I0_9_1_2(op_I0_9_1_2),
    .I0_10_0_0(op_I0_10_0_0),
    .I0_10_0_1(op_I0_10_0_1),
    .I0_10_0_2(op_I0_10_0_2),
    .I0_10_1_0(op_I0_10_1_0),
    .I0_10_1_1(op_I0_10_1_1),
    .I0_10_1_2(op_I0_10_1_2),
    .I0_11_0_0(op_I0_11_0_0),
    .I0_11_0_1(op_I0_11_0_1),
    .I0_11_0_2(op_I0_11_0_2),
    .I0_11_1_0(op_I0_11_1_0),
    .I0_11_1_1(op_I0_11_1_1),
    .I0_11_1_2(op_I0_11_1_2),
    .I0_12_0_0(op_I0_12_0_0),
    .I0_12_0_1(op_I0_12_0_1),
    .I0_12_0_2(op_I0_12_0_2),
    .I0_12_1_0(op_I0_12_1_0),
    .I0_12_1_1(op_I0_12_1_1),
    .I0_12_1_2(op_I0_12_1_2),
    .I0_13_0_0(op_I0_13_0_0),
    .I0_13_0_1(op_I0_13_0_1),
    .I0_13_0_2(op_I0_13_0_2),
    .I0_13_1_0(op_I0_13_1_0),
    .I0_13_1_1(op_I0_13_1_1),
    .I0_13_1_2(op_I0_13_1_2),
    .I0_14_0_0(op_I0_14_0_0),
    .I0_14_0_1(op_I0_14_0_1),
    .I0_14_0_2(op_I0_14_0_2),
    .I0_14_1_0(op_I0_14_1_0),
    .I0_14_1_1(op_I0_14_1_1),
    .I0_14_1_2(op_I0_14_1_2),
    .I0_15_0_0(op_I0_15_0_0),
    .I0_15_0_1(op_I0_15_0_1),
    .I0_15_0_2(op_I0_15_0_2),
    .I0_15_1_0(op_I0_15_1_0),
    .I0_15_1_1(op_I0_15_1_1),
    .I0_15_1_2(op_I0_15_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .I1_8_0(op_I1_8_0),
    .I1_8_1(op_I1_8_1),
    .I1_8_2(op_I1_8_2),
    .I1_9_0(op_I1_9_0),
    .I1_9_1(op_I1_9_1),
    .I1_9_2(op_I1_9_2),
    .I1_10_0(op_I1_10_0),
    .I1_10_1(op_I1_10_1),
    .I1_10_2(op_I1_10_2),
    .I1_11_0(op_I1_11_0),
    .I1_11_1(op_I1_11_1),
    .I1_11_2(op_I1_11_2),
    .I1_12_0(op_I1_12_0),
    .I1_12_1(op_I1_12_1),
    .I1_12_2(op_I1_12_2),
    .I1_13_0(op_I1_13_0),
    .I1_13_1(op_I1_13_1),
    .I1_13_2(op_I1_13_2),
    .I1_14_0(op_I1_14_0),
    .I1_14_1(op_I1_14_1),
    .I1_14_2(op_I1_14_2),
    .I1_15_0(op_I1_15_0),
    .I1_15_1(op_I1_15_1),
    .I1_15_2(op_I1_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_8_2_0(op_O_8_2_0),
    .O_8_2_1(op_O_8_2_1),
    .O_8_2_2(op_O_8_2_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_9_2_0(op_O_9_2_0),
    .O_9_2_1(op_O_9_2_1),
    .O_9_2_2(op_O_9_2_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_10_2_0(op_O_10_2_0),
    .O_10_2_1(op_O_10_2_1),
    .O_10_2_2(op_O_10_2_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_11_2_0(op_O_11_2_0),
    .O_11_2_1(op_O_11_2_1),
    .O_11_2_2(op_O_11_2_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_12_2_0(op_O_12_2_0),
    .O_12_2_1(op_O_12_2_1),
    .O_12_2_2(op_O_12_2_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_13_2_0(op_O_13_2_0),
    .O_13_2_1(op_O_13_2_1),
    .O_13_2_2(op_O_13_2_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_14_2_0(op_O_14_2_0),
    .O_14_2_1(op_O_14_2_1),
    .O_14_2_2(op_O_14_2_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2),
    .O_15_2_0(op_O_15_2_0),
    .O_15_2_1(op_O_15_2_1),
    .O_15_2_2(op_O_15_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_2_0 = op_O_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_2_1 = op_O_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_2_2 = op_O_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_1_2_0 = op_O_1_2_0; // @[Map2T.scala 17:7]
  assign O_1_2_1 = op_O_1_2_1; // @[Map2T.scala 17:7]
  assign O_1_2_2 = op_O_1_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_2_2_0 = op_O_2_2_0; // @[Map2T.scala 17:7]
  assign O_2_2_1 = op_O_2_2_1; // @[Map2T.scala 17:7]
  assign O_2_2_2 = op_O_2_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_3_2_0 = op_O_3_2_0; // @[Map2T.scala 17:7]
  assign O_3_2_1 = op_O_3_2_1; // @[Map2T.scala 17:7]
  assign O_3_2_2 = op_O_3_2_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_4_2_0 = op_O_4_2_0; // @[Map2T.scala 17:7]
  assign O_4_2_1 = op_O_4_2_1; // @[Map2T.scala 17:7]
  assign O_4_2_2 = op_O_4_2_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_5_2_0 = op_O_5_2_0; // @[Map2T.scala 17:7]
  assign O_5_2_1 = op_O_5_2_1; // @[Map2T.scala 17:7]
  assign O_5_2_2 = op_O_5_2_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_6_2_0 = op_O_6_2_0; // @[Map2T.scala 17:7]
  assign O_6_2_1 = op_O_6_2_1; // @[Map2T.scala 17:7]
  assign O_6_2_2 = op_O_6_2_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_7_2_0 = op_O_7_2_0; // @[Map2T.scala 17:7]
  assign O_7_2_1 = op_O_7_2_1; // @[Map2T.scala 17:7]
  assign O_7_2_2 = op_O_7_2_2; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_1 = op_O_8_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_2 = op_O_8_0_2; // @[Map2T.scala 17:7]
  assign O_8_1_0 = op_O_8_1_0; // @[Map2T.scala 17:7]
  assign O_8_1_1 = op_O_8_1_1; // @[Map2T.scala 17:7]
  assign O_8_1_2 = op_O_8_1_2; // @[Map2T.scala 17:7]
  assign O_8_2_0 = op_O_8_2_0; // @[Map2T.scala 17:7]
  assign O_8_2_1 = op_O_8_2_1; // @[Map2T.scala 17:7]
  assign O_8_2_2 = op_O_8_2_2; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_1 = op_O_9_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_2 = op_O_9_0_2; // @[Map2T.scala 17:7]
  assign O_9_1_0 = op_O_9_1_0; // @[Map2T.scala 17:7]
  assign O_9_1_1 = op_O_9_1_1; // @[Map2T.scala 17:7]
  assign O_9_1_2 = op_O_9_1_2; // @[Map2T.scala 17:7]
  assign O_9_2_0 = op_O_9_2_0; // @[Map2T.scala 17:7]
  assign O_9_2_1 = op_O_9_2_1; // @[Map2T.scala 17:7]
  assign O_9_2_2 = op_O_9_2_2; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_1 = op_O_10_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_2 = op_O_10_0_2; // @[Map2T.scala 17:7]
  assign O_10_1_0 = op_O_10_1_0; // @[Map2T.scala 17:7]
  assign O_10_1_1 = op_O_10_1_1; // @[Map2T.scala 17:7]
  assign O_10_1_2 = op_O_10_1_2; // @[Map2T.scala 17:7]
  assign O_10_2_0 = op_O_10_2_0; // @[Map2T.scala 17:7]
  assign O_10_2_1 = op_O_10_2_1; // @[Map2T.scala 17:7]
  assign O_10_2_2 = op_O_10_2_2; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_1 = op_O_11_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_2 = op_O_11_0_2; // @[Map2T.scala 17:7]
  assign O_11_1_0 = op_O_11_1_0; // @[Map2T.scala 17:7]
  assign O_11_1_1 = op_O_11_1_1; // @[Map2T.scala 17:7]
  assign O_11_1_2 = op_O_11_1_2; // @[Map2T.scala 17:7]
  assign O_11_2_0 = op_O_11_2_0; // @[Map2T.scala 17:7]
  assign O_11_2_1 = op_O_11_2_1; // @[Map2T.scala 17:7]
  assign O_11_2_2 = op_O_11_2_2; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_1 = op_O_12_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_2 = op_O_12_0_2; // @[Map2T.scala 17:7]
  assign O_12_1_0 = op_O_12_1_0; // @[Map2T.scala 17:7]
  assign O_12_1_1 = op_O_12_1_1; // @[Map2T.scala 17:7]
  assign O_12_1_2 = op_O_12_1_2; // @[Map2T.scala 17:7]
  assign O_12_2_0 = op_O_12_2_0; // @[Map2T.scala 17:7]
  assign O_12_2_1 = op_O_12_2_1; // @[Map2T.scala 17:7]
  assign O_12_2_2 = op_O_12_2_2; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_1 = op_O_13_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_2 = op_O_13_0_2; // @[Map2T.scala 17:7]
  assign O_13_1_0 = op_O_13_1_0; // @[Map2T.scala 17:7]
  assign O_13_1_1 = op_O_13_1_1; // @[Map2T.scala 17:7]
  assign O_13_1_2 = op_O_13_1_2; // @[Map2T.scala 17:7]
  assign O_13_2_0 = op_O_13_2_0; // @[Map2T.scala 17:7]
  assign O_13_2_1 = op_O_13_2_1; // @[Map2T.scala 17:7]
  assign O_13_2_2 = op_O_13_2_2; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_1 = op_O_14_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_2 = op_O_14_0_2; // @[Map2T.scala 17:7]
  assign O_14_1_0 = op_O_14_1_0; // @[Map2T.scala 17:7]
  assign O_14_1_1 = op_O_14_1_1; // @[Map2T.scala 17:7]
  assign O_14_1_2 = op_O_14_1_2; // @[Map2T.scala 17:7]
  assign O_14_2_0 = op_O_14_2_0; // @[Map2T.scala 17:7]
  assign O_14_2_1 = op_O_14_2_1; // @[Map2T.scala 17:7]
  assign O_14_2_2 = op_O_14_2_2; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_1 = op_O_15_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_2 = op_O_15_0_2; // @[Map2T.scala 17:7]
  assign O_15_1_0 = op_O_15_1_0; // @[Map2T.scala 17:7]
  assign O_15_1_1 = op_O_15_1_1; // @[Map2T.scala 17:7]
  assign O_15_1_2 = op_O_15_1_2; // @[Map2T.scala 17:7]
  assign O_15_2_0 = op_O_15_2_0; // @[Map2T.scala 17:7]
  assign O_15_2_1 = op_O_15_2_1; // @[Map2T.scala 17:7]
  assign O_15_2_2 = op_O_15_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_1_0 = I0_4_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1_1 = I0_4_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_1_2 = I0_4_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_1_0 = I0_5_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1_1 = I0_5_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_1_2 = I0_5_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_1_0 = I0_6_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1_1 = I0_6_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_1_2 = I0_6_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_1_0 = I0_7_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1_1 = I0_7_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_1_2 = I0_7_1_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0 = I0_8_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1 = I0_8_0_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_2 = I0_8_0_2; // @[Map2T.scala 15:11]
  assign op_I0_8_1_0 = I0_8_1_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1_1 = I0_8_1_1; // @[Map2T.scala 15:11]
  assign op_I0_8_1_2 = I0_8_1_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0 = I0_9_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1 = I0_9_0_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_2 = I0_9_0_2; // @[Map2T.scala 15:11]
  assign op_I0_9_1_0 = I0_9_1_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1_1 = I0_9_1_1; // @[Map2T.scala 15:11]
  assign op_I0_9_1_2 = I0_9_1_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0 = I0_10_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1 = I0_10_0_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_2 = I0_10_0_2; // @[Map2T.scala 15:11]
  assign op_I0_10_1_0 = I0_10_1_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1_1 = I0_10_1_1; // @[Map2T.scala 15:11]
  assign op_I0_10_1_2 = I0_10_1_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0 = I0_11_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1 = I0_11_0_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_2 = I0_11_0_2; // @[Map2T.scala 15:11]
  assign op_I0_11_1_0 = I0_11_1_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1_1 = I0_11_1_1; // @[Map2T.scala 15:11]
  assign op_I0_11_1_2 = I0_11_1_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0 = I0_12_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1 = I0_12_0_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_2 = I0_12_0_2; // @[Map2T.scala 15:11]
  assign op_I0_12_1_0 = I0_12_1_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1_1 = I0_12_1_1; // @[Map2T.scala 15:11]
  assign op_I0_12_1_2 = I0_12_1_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0 = I0_13_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1 = I0_13_0_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_2 = I0_13_0_2; // @[Map2T.scala 15:11]
  assign op_I0_13_1_0 = I0_13_1_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1_1 = I0_13_1_1; // @[Map2T.scala 15:11]
  assign op_I0_13_1_2 = I0_13_1_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0 = I0_14_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1 = I0_14_0_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_2 = I0_14_0_2; // @[Map2T.scala 15:11]
  assign op_I0_14_1_0 = I0_14_1_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1_1 = I0_14_1_1; // @[Map2T.scala 15:11]
  assign op_I0_14_1_2 = I0_14_1_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0 = I0_15_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1 = I0_15_0_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_2 = I0_15_0_2; // @[Map2T.scala 15:11]
  assign op_I0_15_1_0 = I0_15_1_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1_1 = I0_15_1_1; // @[Map2T.scala 15:11]
  assign op_I0_15_1_2 = I0_15_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0 = I1_8_0; // @[Map2T.scala 16:11]
  assign op_I1_8_1 = I1_8_1; // @[Map2T.scala 16:11]
  assign op_I1_8_2 = I1_8_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0 = I1_9_0; // @[Map2T.scala 16:11]
  assign op_I1_9_1 = I1_9_1; // @[Map2T.scala 16:11]
  assign op_I1_9_2 = I1_9_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0 = I1_10_0; // @[Map2T.scala 16:11]
  assign op_I1_10_1 = I1_10_1; // @[Map2T.scala 16:11]
  assign op_I1_10_2 = I1_10_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0 = I1_11_0; // @[Map2T.scala 16:11]
  assign op_I1_11_1 = I1_11_1; // @[Map2T.scala 16:11]
  assign op_I1_11_2 = I1_11_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0 = I1_12_0; // @[Map2T.scala 16:11]
  assign op_I1_12_1 = I1_12_1; // @[Map2T.scala 16:11]
  assign op_I1_12_2 = I1_12_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0 = I1_13_0; // @[Map2T.scala 16:11]
  assign op_I1_13_1 = I1_13_1; // @[Map2T.scala 16:11]
  assign op_I1_13_2 = I1_13_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0 = I1_14_0; // @[Map2T.scala 16:11]
  assign op_I1_14_1 = I1_14_1; // @[Map2T.scala 16:11]
  assign op_I1_14_2 = I1_14_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0 = I1_15_0; // @[Map2T.scala 16:11]
  assign op_I1_15_1 = I1_15_1; // @[Map2T.scala 16:11]
  assign op_I1_15_2 = I1_15_2; // @[Map2T.scala 16:11]
endmodule
module PartitionS_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  input  [15:0] I_8_0_0,
  input  [15:0] I_8_0_1,
  input  [15:0] I_8_0_2,
  input  [15:0] I_8_1_0,
  input  [15:0] I_8_1_1,
  input  [15:0] I_8_1_2,
  input  [15:0] I_8_2_0,
  input  [15:0] I_8_2_1,
  input  [15:0] I_8_2_2,
  input  [15:0] I_9_0_0,
  input  [15:0] I_9_0_1,
  input  [15:0] I_9_0_2,
  input  [15:0] I_9_1_0,
  input  [15:0] I_9_1_1,
  input  [15:0] I_9_1_2,
  input  [15:0] I_9_2_0,
  input  [15:0] I_9_2_1,
  input  [15:0] I_9_2_2,
  input  [15:0] I_10_0_0,
  input  [15:0] I_10_0_1,
  input  [15:0] I_10_0_2,
  input  [15:0] I_10_1_0,
  input  [15:0] I_10_1_1,
  input  [15:0] I_10_1_2,
  input  [15:0] I_10_2_0,
  input  [15:0] I_10_2_1,
  input  [15:0] I_10_2_2,
  input  [15:0] I_11_0_0,
  input  [15:0] I_11_0_1,
  input  [15:0] I_11_0_2,
  input  [15:0] I_11_1_0,
  input  [15:0] I_11_1_1,
  input  [15:0] I_11_1_2,
  input  [15:0] I_11_2_0,
  input  [15:0] I_11_2_1,
  input  [15:0] I_11_2_2,
  input  [15:0] I_12_0_0,
  input  [15:0] I_12_0_1,
  input  [15:0] I_12_0_2,
  input  [15:0] I_12_1_0,
  input  [15:0] I_12_1_1,
  input  [15:0] I_12_1_2,
  input  [15:0] I_12_2_0,
  input  [15:0] I_12_2_1,
  input  [15:0] I_12_2_2,
  input  [15:0] I_13_0_0,
  input  [15:0] I_13_0_1,
  input  [15:0] I_13_0_2,
  input  [15:0] I_13_1_0,
  input  [15:0] I_13_1_1,
  input  [15:0] I_13_1_2,
  input  [15:0] I_13_2_0,
  input  [15:0] I_13_2_1,
  input  [15:0] I_13_2_2,
  input  [15:0] I_14_0_0,
  input  [15:0] I_14_0_1,
  input  [15:0] I_14_0_2,
  input  [15:0] I_14_1_0,
  input  [15:0] I_14_1_1,
  input  [15:0] I_14_1_2,
  input  [15:0] I_14_2_0,
  input  [15:0] I_14_2_1,
  input  [15:0] I_14_2_2,
  input  [15:0] I_15_0_0,
  input  [15:0] I_15_0_1,
  input  [15:0] I_15_0_2,
  input  [15:0] I_15_1_0,
  input  [15:0] I_15_1_1,
  input  [15:0] I_15_1_2,
  input  [15:0] I_15_2_0,
  input  [15:0] I_15_2_1,
  input  [15:0] I_15_2_2,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_0_2,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_0_0_1_2,
  output [15:0] O_0_0_2_0,
  output [15:0] O_0_0_2_1,
  output [15:0] O_0_0_2_2,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_0_2,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_1_0_1_2,
  output [15:0] O_1_0_2_0,
  output [15:0] O_1_0_2_1,
  output [15:0] O_1_0_2_2,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_0_2,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_2_0_1_2,
  output [15:0] O_2_0_2_0,
  output [15:0] O_2_0_2_1,
  output [15:0] O_2_0_2_2,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_0_2,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1,
  output [15:0] O_3_0_1_2,
  output [15:0] O_3_0_2_0,
  output [15:0] O_3_0_2_1,
  output [15:0] O_3_0_2_2,
  output [15:0] O_4_0_0_0,
  output [15:0] O_4_0_0_1,
  output [15:0] O_4_0_0_2,
  output [15:0] O_4_0_1_0,
  output [15:0] O_4_0_1_1,
  output [15:0] O_4_0_1_2,
  output [15:0] O_4_0_2_0,
  output [15:0] O_4_0_2_1,
  output [15:0] O_4_0_2_2,
  output [15:0] O_5_0_0_0,
  output [15:0] O_5_0_0_1,
  output [15:0] O_5_0_0_2,
  output [15:0] O_5_0_1_0,
  output [15:0] O_5_0_1_1,
  output [15:0] O_5_0_1_2,
  output [15:0] O_5_0_2_0,
  output [15:0] O_5_0_2_1,
  output [15:0] O_5_0_2_2,
  output [15:0] O_6_0_0_0,
  output [15:0] O_6_0_0_1,
  output [15:0] O_6_0_0_2,
  output [15:0] O_6_0_1_0,
  output [15:0] O_6_0_1_1,
  output [15:0] O_6_0_1_2,
  output [15:0] O_6_0_2_0,
  output [15:0] O_6_0_2_1,
  output [15:0] O_6_0_2_2,
  output [15:0] O_7_0_0_0,
  output [15:0] O_7_0_0_1,
  output [15:0] O_7_0_0_2,
  output [15:0] O_7_0_1_0,
  output [15:0] O_7_0_1_1,
  output [15:0] O_7_0_1_2,
  output [15:0] O_7_0_2_0,
  output [15:0] O_7_0_2_1,
  output [15:0] O_7_0_2_2,
  output [15:0] O_8_0_0_0,
  output [15:0] O_8_0_0_1,
  output [15:0] O_8_0_0_2,
  output [15:0] O_8_0_1_0,
  output [15:0] O_8_0_1_1,
  output [15:0] O_8_0_1_2,
  output [15:0] O_8_0_2_0,
  output [15:0] O_8_0_2_1,
  output [15:0] O_8_0_2_2,
  output [15:0] O_9_0_0_0,
  output [15:0] O_9_0_0_1,
  output [15:0] O_9_0_0_2,
  output [15:0] O_9_0_1_0,
  output [15:0] O_9_0_1_1,
  output [15:0] O_9_0_1_2,
  output [15:0] O_9_0_2_0,
  output [15:0] O_9_0_2_1,
  output [15:0] O_9_0_2_2,
  output [15:0] O_10_0_0_0,
  output [15:0] O_10_0_0_1,
  output [15:0] O_10_0_0_2,
  output [15:0] O_10_0_1_0,
  output [15:0] O_10_0_1_1,
  output [15:0] O_10_0_1_2,
  output [15:0] O_10_0_2_0,
  output [15:0] O_10_0_2_1,
  output [15:0] O_10_0_2_2,
  output [15:0] O_11_0_0_0,
  output [15:0] O_11_0_0_1,
  output [15:0] O_11_0_0_2,
  output [15:0] O_11_0_1_0,
  output [15:0] O_11_0_1_1,
  output [15:0] O_11_0_1_2,
  output [15:0] O_11_0_2_0,
  output [15:0] O_11_0_2_1,
  output [15:0] O_11_0_2_2,
  output [15:0] O_12_0_0_0,
  output [15:0] O_12_0_0_1,
  output [15:0] O_12_0_0_2,
  output [15:0] O_12_0_1_0,
  output [15:0] O_12_0_1_1,
  output [15:0] O_12_0_1_2,
  output [15:0] O_12_0_2_0,
  output [15:0] O_12_0_2_1,
  output [15:0] O_12_0_2_2,
  output [15:0] O_13_0_0_0,
  output [15:0] O_13_0_0_1,
  output [15:0] O_13_0_0_2,
  output [15:0] O_13_0_1_0,
  output [15:0] O_13_0_1_1,
  output [15:0] O_13_0_1_2,
  output [15:0] O_13_0_2_0,
  output [15:0] O_13_0_2_1,
  output [15:0] O_13_0_2_2,
  output [15:0] O_14_0_0_0,
  output [15:0] O_14_0_0_1,
  output [15:0] O_14_0_0_2,
  output [15:0] O_14_0_1_0,
  output [15:0] O_14_0_1_1,
  output [15:0] O_14_0_1_2,
  output [15:0] O_14_0_2_0,
  output [15:0] O_14_0_2_1,
  output [15:0] O_14_0_2_2,
  output [15:0] O_15_0_0_0,
  output [15:0] O_15_0_0_1,
  output [15:0] O_15_0_0_2,
  output [15:0] O_15_0_1_0,
  output [15:0] O_15_0_1_1,
  output [15:0] O_15_0_1_2,
  output [15:0] O_15_0_2_0,
  output [15:0] O_15_0_2_1,
  output [15:0] O_15_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_0_2 = I_2_0_2; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_2_0_1_2 = I_2_1_2; // @[Partition.scala 15:39]
  assign O_2_0_2_0 = I_2_2_0; // @[Partition.scala 15:39]
  assign O_2_0_2_1 = I_2_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2_2 = I_2_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_0_2 = I_3_0_2; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_3_0_1_2 = I_3_1_2; // @[Partition.scala 15:39]
  assign O_3_0_2_0 = I_3_2_0; // @[Partition.scala 15:39]
  assign O_3_0_2_1 = I_3_2_1; // @[Partition.scala 15:39]
  assign O_3_0_2_2 = I_3_2_2; // @[Partition.scala 15:39]
  assign O_4_0_0_0 = I_4_0_0; // @[Partition.scala 15:39]
  assign O_4_0_0_1 = I_4_0_1; // @[Partition.scala 15:39]
  assign O_4_0_0_2 = I_4_0_2; // @[Partition.scala 15:39]
  assign O_4_0_1_0 = I_4_1_0; // @[Partition.scala 15:39]
  assign O_4_0_1_1 = I_4_1_1; // @[Partition.scala 15:39]
  assign O_4_0_1_2 = I_4_1_2; // @[Partition.scala 15:39]
  assign O_4_0_2_0 = I_4_2_0; // @[Partition.scala 15:39]
  assign O_4_0_2_1 = I_4_2_1; // @[Partition.scala 15:39]
  assign O_4_0_2_2 = I_4_2_2; // @[Partition.scala 15:39]
  assign O_5_0_0_0 = I_5_0_0; // @[Partition.scala 15:39]
  assign O_5_0_0_1 = I_5_0_1; // @[Partition.scala 15:39]
  assign O_5_0_0_2 = I_5_0_2; // @[Partition.scala 15:39]
  assign O_5_0_1_0 = I_5_1_0; // @[Partition.scala 15:39]
  assign O_5_0_1_1 = I_5_1_1; // @[Partition.scala 15:39]
  assign O_5_0_1_2 = I_5_1_2; // @[Partition.scala 15:39]
  assign O_5_0_2_0 = I_5_2_0; // @[Partition.scala 15:39]
  assign O_5_0_2_1 = I_5_2_1; // @[Partition.scala 15:39]
  assign O_5_0_2_2 = I_5_2_2; // @[Partition.scala 15:39]
  assign O_6_0_0_0 = I_6_0_0; // @[Partition.scala 15:39]
  assign O_6_0_0_1 = I_6_0_1; // @[Partition.scala 15:39]
  assign O_6_0_0_2 = I_6_0_2; // @[Partition.scala 15:39]
  assign O_6_0_1_0 = I_6_1_0; // @[Partition.scala 15:39]
  assign O_6_0_1_1 = I_6_1_1; // @[Partition.scala 15:39]
  assign O_6_0_1_2 = I_6_1_2; // @[Partition.scala 15:39]
  assign O_6_0_2_0 = I_6_2_0; // @[Partition.scala 15:39]
  assign O_6_0_2_1 = I_6_2_1; // @[Partition.scala 15:39]
  assign O_6_0_2_2 = I_6_2_2; // @[Partition.scala 15:39]
  assign O_7_0_0_0 = I_7_0_0; // @[Partition.scala 15:39]
  assign O_7_0_0_1 = I_7_0_1; // @[Partition.scala 15:39]
  assign O_7_0_0_2 = I_7_0_2; // @[Partition.scala 15:39]
  assign O_7_0_1_0 = I_7_1_0; // @[Partition.scala 15:39]
  assign O_7_0_1_1 = I_7_1_1; // @[Partition.scala 15:39]
  assign O_7_0_1_2 = I_7_1_2; // @[Partition.scala 15:39]
  assign O_7_0_2_0 = I_7_2_0; // @[Partition.scala 15:39]
  assign O_7_0_2_1 = I_7_2_1; // @[Partition.scala 15:39]
  assign O_7_0_2_2 = I_7_2_2; // @[Partition.scala 15:39]
  assign O_8_0_0_0 = I_8_0_0; // @[Partition.scala 15:39]
  assign O_8_0_0_1 = I_8_0_1; // @[Partition.scala 15:39]
  assign O_8_0_0_2 = I_8_0_2; // @[Partition.scala 15:39]
  assign O_8_0_1_0 = I_8_1_0; // @[Partition.scala 15:39]
  assign O_8_0_1_1 = I_8_1_1; // @[Partition.scala 15:39]
  assign O_8_0_1_2 = I_8_1_2; // @[Partition.scala 15:39]
  assign O_8_0_2_0 = I_8_2_0; // @[Partition.scala 15:39]
  assign O_8_0_2_1 = I_8_2_1; // @[Partition.scala 15:39]
  assign O_8_0_2_2 = I_8_2_2; // @[Partition.scala 15:39]
  assign O_9_0_0_0 = I_9_0_0; // @[Partition.scala 15:39]
  assign O_9_0_0_1 = I_9_0_1; // @[Partition.scala 15:39]
  assign O_9_0_0_2 = I_9_0_2; // @[Partition.scala 15:39]
  assign O_9_0_1_0 = I_9_1_0; // @[Partition.scala 15:39]
  assign O_9_0_1_1 = I_9_1_1; // @[Partition.scala 15:39]
  assign O_9_0_1_2 = I_9_1_2; // @[Partition.scala 15:39]
  assign O_9_0_2_0 = I_9_2_0; // @[Partition.scala 15:39]
  assign O_9_0_2_1 = I_9_2_1; // @[Partition.scala 15:39]
  assign O_9_0_2_2 = I_9_2_2; // @[Partition.scala 15:39]
  assign O_10_0_0_0 = I_10_0_0; // @[Partition.scala 15:39]
  assign O_10_0_0_1 = I_10_0_1; // @[Partition.scala 15:39]
  assign O_10_0_0_2 = I_10_0_2; // @[Partition.scala 15:39]
  assign O_10_0_1_0 = I_10_1_0; // @[Partition.scala 15:39]
  assign O_10_0_1_1 = I_10_1_1; // @[Partition.scala 15:39]
  assign O_10_0_1_2 = I_10_1_2; // @[Partition.scala 15:39]
  assign O_10_0_2_0 = I_10_2_0; // @[Partition.scala 15:39]
  assign O_10_0_2_1 = I_10_2_1; // @[Partition.scala 15:39]
  assign O_10_0_2_2 = I_10_2_2; // @[Partition.scala 15:39]
  assign O_11_0_0_0 = I_11_0_0; // @[Partition.scala 15:39]
  assign O_11_0_0_1 = I_11_0_1; // @[Partition.scala 15:39]
  assign O_11_0_0_2 = I_11_0_2; // @[Partition.scala 15:39]
  assign O_11_0_1_0 = I_11_1_0; // @[Partition.scala 15:39]
  assign O_11_0_1_1 = I_11_1_1; // @[Partition.scala 15:39]
  assign O_11_0_1_2 = I_11_1_2; // @[Partition.scala 15:39]
  assign O_11_0_2_0 = I_11_2_0; // @[Partition.scala 15:39]
  assign O_11_0_2_1 = I_11_2_1; // @[Partition.scala 15:39]
  assign O_11_0_2_2 = I_11_2_2; // @[Partition.scala 15:39]
  assign O_12_0_0_0 = I_12_0_0; // @[Partition.scala 15:39]
  assign O_12_0_0_1 = I_12_0_1; // @[Partition.scala 15:39]
  assign O_12_0_0_2 = I_12_0_2; // @[Partition.scala 15:39]
  assign O_12_0_1_0 = I_12_1_0; // @[Partition.scala 15:39]
  assign O_12_0_1_1 = I_12_1_1; // @[Partition.scala 15:39]
  assign O_12_0_1_2 = I_12_1_2; // @[Partition.scala 15:39]
  assign O_12_0_2_0 = I_12_2_0; // @[Partition.scala 15:39]
  assign O_12_0_2_1 = I_12_2_1; // @[Partition.scala 15:39]
  assign O_12_0_2_2 = I_12_2_2; // @[Partition.scala 15:39]
  assign O_13_0_0_0 = I_13_0_0; // @[Partition.scala 15:39]
  assign O_13_0_0_1 = I_13_0_1; // @[Partition.scala 15:39]
  assign O_13_0_0_2 = I_13_0_2; // @[Partition.scala 15:39]
  assign O_13_0_1_0 = I_13_1_0; // @[Partition.scala 15:39]
  assign O_13_0_1_1 = I_13_1_1; // @[Partition.scala 15:39]
  assign O_13_0_1_2 = I_13_1_2; // @[Partition.scala 15:39]
  assign O_13_0_2_0 = I_13_2_0; // @[Partition.scala 15:39]
  assign O_13_0_2_1 = I_13_2_1; // @[Partition.scala 15:39]
  assign O_13_0_2_2 = I_13_2_2; // @[Partition.scala 15:39]
  assign O_14_0_0_0 = I_14_0_0; // @[Partition.scala 15:39]
  assign O_14_0_0_1 = I_14_0_1; // @[Partition.scala 15:39]
  assign O_14_0_0_2 = I_14_0_2; // @[Partition.scala 15:39]
  assign O_14_0_1_0 = I_14_1_0; // @[Partition.scala 15:39]
  assign O_14_0_1_1 = I_14_1_1; // @[Partition.scala 15:39]
  assign O_14_0_1_2 = I_14_1_2; // @[Partition.scala 15:39]
  assign O_14_0_2_0 = I_14_2_0; // @[Partition.scala 15:39]
  assign O_14_0_2_1 = I_14_2_1; // @[Partition.scala 15:39]
  assign O_14_0_2_2 = I_14_2_2; // @[Partition.scala 15:39]
  assign O_15_0_0_0 = I_15_0_0; // @[Partition.scala 15:39]
  assign O_15_0_0_1 = I_15_0_1; // @[Partition.scala 15:39]
  assign O_15_0_0_2 = I_15_0_2; // @[Partition.scala 15:39]
  assign O_15_0_1_0 = I_15_1_0; // @[Partition.scala 15:39]
  assign O_15_0_1_1 = I_15_1_1; // @[Partition.scala 15:39]
  assign O_15_0_1_2 = I_15_1_2; // @[Partition.scala 15:39]
  assign O_15_0_2_0 = I_15_2_0; // @[Partition.scala 15:39]
  assign O_15_0_2_1 = I_15_2_1; // @[Partition.scala 15:39]
  assign O_15_0_2_2 = I_15_2_2; // @[Partition.scala 15:39]
endmodule
module MapT_6(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  input  [15:0] I_8_0_0,
  input  [15:0] I_8_0_1,
  input  [15:0] I_8_0_2,
  input  [15:0] I_8_1_0,
  input  [15:0] I_8_1_1,
  input  [15:0] I_8_1_2,
  input  [15:0] I_8_2_0,
  input  [15:0] I_8_2_1,
  input  [15:0] I_8_2_2,
  input  [15:0] I_9_0_0,
  input  [15:0] I_9_0_1,
  input  [15:0] I_9_0_2,
  input  [15:0] I_9_1_0,
  input  [15:0] I_9_1_1,
  input  [15:0] I_9_1_2,
  input  [15:0] I_9_2_0,
  input  [15:0] I_9_2_1,
  input  [15:0] I_9_2_2,
  input  [15:0] I_10_0_0,
  input  [15:0] I_10_0_1,
  input  [15:0] I_10_0_2,
  input  [15:0] I_10_1_0,
  input  [15:0] I_10_1_1,
  input  [15:0] I_10_1_2,
  input  [15:0] I_10_2_0,
  input  [15:0] I_10_2_1,
  input  [15:0] I_10_2_2,
  input  [15:0] I_11_0_0,
  input  [15:0] I_11_0_1,
  input  [15:0] I_11_0_2,
  input  [15:0] I_11_1_0,
  input  [15:0] I_11_1_1,
  input  [15:0] I_11_1_2,
  input  [15:0] I_11_2_0,
  input  [15:0] I_11_2_1,
  input  [15:0] I_11_2_2,
  input  [15:0] I_12_0_0,
  input  [15:0] I_12_0_1,
  input  [15:0] I_12_0_2,
  input  [15:0] I_12_1_0,
  input  [15:0] I_12_1_1,
  input  [15:0] I_12_1_2,
  input  [15:0] I_12_2_0,
  input  [15:0] I_12_2_1,
  input  [15:0] I_12_2_2,
  input  [15:0] I_13_0_0,
  input  [15:0] I_13_0_1,
  input  [15:0] I_13_0_2,
  input  [15:0] I_13_1_0,
  input  [15:0] I_13_1_1,
  input  [15:0] I_13_1_2,
  input  [15:0] I_13_2_0,
  input  [15:0] I_13_2_1,
  input  [15:0] I_13_2_2,
  input  [15:0] I_14_0_0,
  input  [15:0] I_14_0_1,
  input  [15:0] I_14_0_2,
  input  [15:0] I_14_1_0,
  input  [15:0] I_14_1_1,
  input  [15:0] I_14_1_2,
  input  [15:0] I_14_2_0,
  input  [15:0] I_14_2_1,
  input  [15:0] I_14_2_2,
  input  [15:0] I_15_0_0,
  input  [15:0] I_15_0_1,
  input  [15:0] I_15_0_2,
  input  [15:0] I_15_1_0,
  input  [15:0] I_15_1_1,
  input  [15:0] I_15_1_2,
  input  [15:0] I_15_2_0,
  input  [15:0] I_15_2_1,
  input  [15:0] I_15_2_2,
  output [15:0] O_0_0_0_0,
  output [15:0] O_0_0_0_1,
  output [15:0] O_0_0_0_2,
  output [15:0] O_0_0_1_0,
  output [15:0] O_0_0_1_1,
  output [15:0] O_0_0_1_2,
  output [15:0] O_0_0_2_0,
  output [15:0] O_0_0_2_1,
  output [15:0] O_0_0_2_2,
  output [15:0] O_1_0_0_0,
  output [15:0] O_1_0_0_1,
  output [15:0] O_1_0_0_2,
  output [15:0] O_1_0_1_0,
  output [15:0] O_1_0_1_1,
  output [15:0] O_1_0_1_2,
  output [15:0] O_1_0_2_0,
  output [15:0] O_1_0_2_1,
  output [15:0] O_1_0_2_2,
  output [15:0] O_2_0_0_0,
  output [15:0] O_2_0_0_1,
  output [15:0] O_2_0_0_2,
  output [15:0] O_2_0_1_0,
  output [15:0] O_2_0_1_1,
  output [15:0] O_2_0_1_2,
  output [15:0] O_2_0_2_0,
  output [15:0] O_2_0_2_1,
  output [15:0] O_2_0_2_2,
  output [15:0] O_3_0_0_0,
  output [15:0] O_3_0_0_1,
  output [15:0] O_3_0_0_2,
  output [15:0] O_3_0_1_0,
  output [15:0] O_3_0_1_1,
  output [15:0] O_3_0_1_2,
  output [15:0] O_3_0_2_0,
  output [15:0] O_3_0_2_1,
  output [15:0] O_3_0_2_2,
  output [15:0] O_4_0_0_0,
  output [15:0] O_4_0_0_1,
  output [15:0] O_4_0_0_2,
  output [15:0] O_4_0_1_0,
  output [15:0] O_4_0_1_1,
  output [15:0] O_4_0_1_2,
  output [15:0] O_4_0_2_0,
  output [15:0] O_4_0_2_1,
  output [15:0] O_4_0_2_2,
  output [15:0] O_5_0_0_0,
  output [15:0] O_5_0_0_1,
  output [15:0] O_5_0_0_2,
  output [15:0] O_5_0_1_0,
  output [15:0] O_5_0_1_1,
  output [15:0] O_5_0_1_2,
  output [15:0] O_5_0_2_0,
  output [15:0] O_5_0_2_1,
  output [15:0] O_5_0_2_2,
  output [15:0] O_6_0_0_0,
  output [15:0] O_6_0_0_1,
  output [15:0] O_6_0_0_2,
  output [15:0] O_6_0_1_0,
  output [15:0] O_6_0_1_1,
  output [15:0] O_6_0_1_2,
  output [15:0] O_6_0_2_0,
  output [15:0] O_6_0_2_1,
  output [15:0] O_6_0_2_2,
  output [15:0] O_7_0_0_0,
  output [15:0] O_7_0_0_1,
  output [15:0] O_7_0_0_2,
  output [15:0] O_7_0_1_0,
  output [15:0] O_7_0_1_1,
  output [15:0] O_7_0_1_2,
  output [15:0] O_7_0_2_0,
  output [15:0] O_7_0_2_1,
  output [15:0] O_7_0_2_2,
  output [15:0] O_8_0_0_0,
  output [15:0] O_8_0_0_1,
  output [15:0] O_8_0_0_2,
  output [15:0] O_8_0_1_0,
  output [15:0] O_8_0_1_1,
  output [15:0] O_8_0_1_2,
  output [15:0] O_8_0_2_0,
  output [15:0] O_8_0_2_1,
  output [15:0] O_8_0_2_2,
  output [15:0] O_9_0_0_0,
  output [15:0] O_9_0_0_1,
  output [15:0] O_9_0_0_2,
  output [15:0] O_9_0_1_0,
  output [15:0] O_9_0_1_1,
  output [15:0] O_9_0_1_2,
  output [15:0] O_9_0_2_0,
  output [15:0] O_9_0_2_1,
  output [15:0] O_9_0_2_2,
  output [15:0] O_10_0_0_0,
  output [15:0] O_10_0_0_1,
  output [15:0] O_10_0_0_2,
  output [15:0] O_10_0_1_0,
  output [15:0] O_10_0_1_1,
  output [15:0] O_10_0_1_2,
  output [15:0] O_10_0_2_0,
  output [15:0] O_10_0_2_1,
  output [15:0] O_10_0_2_2,
  output [15:0] O_11_0_0_0,
  output [15:0] O_11_0_0_1,
  output [15:0] O_11_0_0_2,
  output [15:0] O_11_0_1_0,
  output [15:0] O_11_0_1_1,
  output [15:0] O_11_0_1_2,
  output [15:0] O_11_0_2_0,
  output [15:0] O_11_0_2_1,
  output [15:0] O_11_0_2_2,
  output [15:0] O_12_0_0_0,
  output [15:0] O_12_0_0_1,
  output [15:0] O_12_0_0_2,
  output [15:0] O_12_0_1_0,
  output [15:0] O_12_0_1_1,
  output [15:0] O_12_0_1_2,
  output [15:0] O_12_0_2_0,
  output [15:0] O_12_0_2_1,
  output [15:0] O_12_0_2_2,
  output [15:0] O_13_0_0_0,
  output [15:0] O_13_0_0_1,
  output [15:0] O_13_0_0_2,
  output [15:0] O_13_0_1_0,
  output [15:0] O_13_0_1_1,
  output [15:0] O_13_0_1_2,
  output [15:0] O_13_0_2_0,
  output [15:0] O_13_0_2_1,
  output [15:0] O_13_0_2_2,
  output [15:0] O_14_0_0_0,
  output [15:0] O_14_0_0_1,
  output [15:0] O_14_0_0_2,
  output [15:0] O_14_0_1_0,
  output [15:0] O_14_0_1_1,
  output [15:0] O_14_0_1_2,
  output [15:0] O_14_0_2_0,
  output [15:0] O_14_0_2_1,
  output [15:0] O_14_0_2_2,
  output [15:0] O_15_0_0_0,
  output [15:0] O_15_0_0_1,
  output [15:0] O_15_0_0_2,
  output [15:0] O_15_0_1_0,
  output [15:0] O_15_0_1_1,
  output [15:0] O_15_0_1_2,
  output [15:0] O_15_0_2_0,
  output [15:0] O_15_0_2_1,
  output [15:0] O_15_0_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_2_2; // @[MapT.scala 8:20]
  PartitionS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_8_1_2(op_I_8_1_2),
    .I_8_2_0(op_I_8_2_0),
    .I_8_2_1(op_I_8_2_1),
    .I_8_2_2(op_I_8_2_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_9_1_2(op_I_9_1_2),
    .I_9_2_0(op_I_9_2_0),
    .I_9_2_1(op_I_9_2_1),
    .I_9_2_2(op_I_9_2_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_10_1_2(op_I_10_1_2),
    .I_10_2_0(op_I_10_2_0),
    .I_10_2_1(op_I_10_2_1),
    .I_10_2_2(op_I_10_2_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_11_1_2(op_I_11_1_2),
    .I_11_2_0(op_I_11_2_0),
    .I_11_2_1(op_I_11_2_1),
    .I_11_2_2(op_I_11_2_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_12_1_2(op_I_12_1_2),
    .I_12_2_0(op_I_12_2_0),
    .I_12_2_1(op_I_12_2_1),
    .I_12_2_2(op_I_12_2_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_13_1_2(op_I_13_1_2),
    .I_13_2_0(op_I_13_2_0),
    .I_13_2_1(op_I_13_2_1),
    .I_13_2_2(op_I_13_2_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_14_1_2(op_I_14_1_2),
    .I_14_2_0(op_I_14_2_0),
    .I_14_2_1(op_I_14_2_1),
    .I_14_2_2(op_I_14_2_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .I_15_1_2(op_I_15_1_2),
    .I_15_2_0(op_I_15_2_0),
    .I_15_2_1(op_I_15_2_1),
    .I_15_2_2(op_I_15_2_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_4_0_2_0(op_O_4_0_2_0),
    .O_4_0_2_1(op_O_4_0_2_1),
    .O_4_0_2_2(op_O_4_0_2_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_5_0_2_0(op_O_5_0_2_0),
    .O_5_0_2_1(op_O_5_0_2_1),
    .O_5_0_2_2(op_O_5_0_2_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_6_0_2_0(op_O_6_0_2_0),
    .O_6_0_2_1(op_O_6_0_2_1),
    .O_6_0_2_2(op_O_6_0_2_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_7_0_2_0(op_O_7_0_2_0),
    .O_7_0_2_1(op_O_7_0_2_1),
    .O_7_0_2_2(op_O_7_0_2_2),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_8_0_0_2(op_O_8_0_0_2),
    .O_8_0_1_0(op_O_8_0_1_0),
    .O_8_0_1_1(op_O_8_0_1_1),
    .O_8_0_1_2(op_O_8_0_1_2),
    .O_8_0_2_0(op_O_8_0_2_0),
    .O_8_0_2_1(op_O_8_0_2_1),
    .O_8_0_2_2(op_O_8_0_2_2),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_9_0_0_2(op_O_9_0_0_2),
    .O_9_0_1_0(op_O_9_0_1_0),
    .O_9_0_1_1(op_O_9_0_1_1),
    .O_9_0_1_2(op_O_9_0_1_2),
    .O_9_0_2_0(op_O_9_0_2_0),
    .O_9_0_2_1(op_O_9_0_2_1),
    .O_9_0_2_2(op_O_9_0_2_2),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_10_0_0_2(op_O_10_0_0_2),
    .O_10_0_1_0(op_O_10_0_1_0),
    .O_10_0_1_1(op_O_10_0_1_1),
    .O_10_0_1_2(op_O_10_0_1_2),
    .O_10_0_2_0(op_O_10_0_2_0),
    .O_10_0_2_1(op_O_10_0_2_1),
    .O_10_0_2_2(op_O_10_0_2_2),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_11_0_0_2(op_O_11_0_0_2),
    .O_11_0_1_0(op_O_11_0_1_0),
    .O_11_0_1_1(op_O_11_0_1_1),
    .O_11_0_1_2(op_O_11_0_1_2),
    .O_11_0_2_0(op_O_11_0_2_0),
    .O_11_0_2_1(op_O_11_0_2_1),
    .O_11_0_2_2(op_O_11_0_2_2),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_12_0_0_2(op_O_12_0_0_2),
    .O_12_0_1_0(op_O_12_0_1_0),
    .O_12_0_1_1(op_O_12_0_1_1),
    .O_12_0_1_2(op_O_12_0_1_2),
    .O_12_0_2_0(op_O_12_0_2_0),
    .O_12_0_2_1(op_O_12_0_2_1),
    .O_12_0_2_2(op_O_12_0_2_2),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_13_0_0_2(op_O_13_0_0_2),
    .O_13_0_1_0(op_O_13_0_1_0),
    .O_13_0_1_1(op_O_13_0_1_1),
    .O_13_0_1_2(op_O_13_0_1_2),
    .O_13_0_2_0(op_O_13_0_2_0),
    .O_13_0_2_1(op_O_13_0_2_1),
    .O_13_0_2_2(op_O_13_0_2_2),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_14_0_0_2(op_O_14_0_0_2),
    .O_14_0_1_0(op_O_14_0_1_0),
    .O_14_0_1_1(op_O_14_0_1_1),
    .O_14_0_1_2(op_O_14_0_1_2),
    .O_14_0_2_0(op_O_14_0_2_0),
    .O_14_0_2_1(op_O_14_0_2_1),
    .O_14_0_2_2(op_O_14_0_2_2),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1),
    .O_15_0_0_2(op_O_15_0_0_2),
    .O_15_0_1_0(op_O_15_0_1_0),
    .O_15_0_1_1(op_O_15_0_1_1),
    .O_15_0_1_2(op_O_15_0_1_2),
    .O_15_0_2_0(op_O_15_0_2_0),
    .O_15_0_2_1(op_O_15_0_2_1),
    .O_15_0_2_2(op_O_15_0_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[MapT.scala 15:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[MapT.scala 15:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[MapT.scala 15:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[MapT.scala 15:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[MapT.scala 15:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[MapT.scala 15:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[MapT.scala 15:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[MapT.scala 15:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[MapT.scala 15:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[MapT.scala 15:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[MapT.scala 15:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[MapT.scala 15:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[MapT.scala 15:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[MapT.scala 15:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[MapT.scala 15:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[MapT.scala 15:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[MapT.scala 15:7]
  assign O_4_0_2_0 = op_O_4_0_2_0; // @[MapT.scala 15:7]
  assign O_4_0_2_1 = op_O_4_0_2_1; // @[MapT.scala 15:7]
  assign O_4_0_2_2 = op_O_4_0_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[MapT.scala 15:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[MapT.scala 15:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[MapT.scala 15:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[MapT.scala 15:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[MapT.scala 15:7]
  assign O_5_0_2_0 = op_O_5_0_2_0; // @[MapT.scala 15:7]
  assign O_5_0_2_1 = op_O_5_0_2_1; // @[MapT.scala 15:7]
  assign O_5_0_2_2 = op_O_5_0_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[MapT.scala 15:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[MapT.scala 15:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[MapT.scala 15:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[MapT.scala 15:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[MapT.scala 15:7]
  assign O_6_0_2_0 = op_O_6_0_2_0; // @[MapT.scala 15:7]
  assign O_6_0_2_1 = op_O_6_0_2_1; // @[MapT.scala 15:7]
  assign O_6_0_2_2 = op_O_6_0_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[MapT.scala 15:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[MapT.scala 15:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[MapT.scala 15:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[MapT.scala 15:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[MapT.scala 15:7]
  assign O_7_0_2_0 = op_O_7_0_2_0; // @[MapT.scala 15:7]
  assign O_7_0_2_1 = op_O_7_0_2_1; // @[MapT.scala 15:7]
  assign O_7_0_2_2 = op_O_7_0_2_2; // @[MapT.scala 15:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[MapT.scala 15:7]
  assign O_8_0_0_2 = op_O_8_0_0_2; // @[MapT.scala 15:7]
  assign O_8_0_1_0 = op_O_8_0_1_0; // @[MapT.scala 15:7]
  assign O_8_0_1_1 = op_O_8_0_1_1; // @[MapT.scala 15:7]
  assign O_8_0_1_2 = op_O_8_0_1_2; // @[MapT.scala 15:7]
  assign O_8_0_2_0 = op_O_8_0_2_0; // @[MapT.scala 15:7]
  assign O_8_0_2_1 = op_O_8_0_2_1; // @[MapT.scala 15:7]
  assign O_8_0_2_2 = op_O_8_0_2_2; // @[MapT.scala 15:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[MapT.scala 15:7]
  assign O_9_0_0_2 = op_O_9_0_0_2; // @[MapT.scala 15:7]
  assign O_9_0_1_0 = op_O_9_0_1_0; // @[MapT.scala 15:7]
  assign O_9_0_1_1 = op_O_9_0_1_1; // @[MapT.scala 15:7]
  assign O_9_0_1_2 = op_O_9_0_1_2; // @[MapT.scala 15:7]
  assign O_9_0_2_0 = op_O_9_0_2_0; // @[MapT.scala 15:7]
  assign O_9_0_2_1 = op_O_9_0_2_1; // @[MapT.scala 15:7]
  assign O_9_0_2_2 = op_O_9_0_2_2; // @[MapT.scala 15:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[MapT.scala 15:7]
  assign O_10_0_0_2 = op_O_10_0_0_2; // @[MapT.scala 15:7]
  assign O_10_0_1_0 = op_O_10_0_1_0; // @[MapT.scala 15:7]
  assign O_10_0_1_1 = op_O_10_0_1_1; // @[MapT.scala 15:7]
  assign O_10_0_1_2 = op_O_10_0_1_2; // @[MapT.scala 15:7]
  assign O_10_0_2_0 = op_O_10_0_2_0; // @[MapT.scala 15:7]
  assign O_10_0_2_1 = op_O_10_0_2_1; // @[MapT.scala 15:7]
  assign O_10_0_2_2 = op_O_10_0_2_2; // @[MapT.scala 15:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[MapT.scala 15:7]
  assign O_11_0_0_2 = op_O_11_0_0_2; // @[MapT.scala 15:7]
  assign O_11_0_1_0 = op_O_11_0_1_0; // @[MapT.scala 15:7]
  assign O_11_0_1_1 = op_O_11_0_1_1; // @[MapT.scala 15:7]
  assign O_11_0_1_2 = op_O_11_0_1_2; // @[MapT.scala 15:7]
  assign O_11_0_2_0 = op_O_11_0_2_0; // @[MapT.scala 15:7]
  assign O_11_0_2_1 = op_O_11_0_2_1; // @[MapT.scala 15:7]
  assign O_11_0_2_2 = op_O_11_0_2_2; // @[MapT.scala 15:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[MapT.scala 15:7]
  assign O_12_0_0_2 = op_O_12_0_0_2; // @[MapT.scala 15:7]
  assign O_12_0_1_0 = op_O_12_0_1_0; // @[MapT.scala 15:7]
  assign O_12_0_1_1 = op_O_12_0_1_1; // @[MapT.scala 15:7]
  assign O_12_0_1_2 = op_O_12_0_1_2; // @[MapT.scala 15:7]
  assign O_12_0_2_0 = op_O_12_0_2_0; // @[MapT.scala 15:7]
  assign O_12_0_2_1 = op_O_12_0_2_1; // @[MapT.scala 15:7]
  assign O_12_0_2_2 = op_O_12_0_2_2; // @[MapT.scala 15:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[MapT.scala 15:7]
  assign O_13_0_0_2 = op_O_13_0_0_2; // @[MapT.scala 15:7]
  assign O_13_0_1_0 = op_O_13_0_1_0; // @[MapT.scala 15:7]
  assign O_13_0_1_1 = op_O_13_0_1_1; // @[MapT.scala 15:7]
  assign O_13_0_1_2 = op_O_13_0_1_2; // @[MapT.scala 15:7]
  assign O_13_0_2_0 = op_O_13_0_2_0; // @[MapT.scala 15:7]
  assign O_13_0_2_1 = op_O_13_0_2_1; // @[MapT.scala 15:7]
  assign O_13_0_2_2 = op_O_13_0_2_2; // @[MapT.scala 15:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[MapT.scala 15:7]
  assign O_14_0_0_2 = op_O_14_0_0_2; // @[MapT.scala 15:7]
  assign O_14_0_1_0 = op_O_14_0_1_0; // @[MapT.scala 15:7]
  assign O_14_0_1_1 = op_O_14_0_1_1; // @[MapT.scala 15:7]
  assign O_14_0_1_2 = op_O_14_0_1_2; // @[MapT.scala 15:7]
  assign O_14_0_2_0 = op_O_14_0_2_0; // @[MapT.scala 15:7]
  assign O_14_0_2_1 = op_O_14_0_2_1; // @[MapT.scala 15:7]
  assign O_14_0_2_2 = op_O_14_0_2_2; // @[MapT.scala 15:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[MapT.scala 15:7]
  assign O_15_0_0_2 = op_O_15_0_0_2; // @[MapT.scala 15:7]
  assign O_15_0_1_0 = op_O_15_0_1_0; // @[MapT.scala 15:7]
  assign O_15_0_1_1 = op_O_15_0_1_1; // @[MapT.scala 15:7]
  assign O_15_0_1_2 = op_O_15_0_1_2; // @[MapT.scala 15:7]
  assign O_15_0_2_0 = op_O_15_0_2_0; // @[MapT.scala 15:7]
  assign O_15_0_2_1 = op_O_15_0_2_1; // @[MapT.scala 15:7]
  assign O_15_0_2_2 = op_O_15_0_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_8_1_2 = I_8_1_2; // @[MapT.scala 14:10]
  assign op_I_8_2_0 = I_8_2_0; // @[MapT.scala 14:10]
  assign op_I_8_2_1 = I_8_2_1; // @[MapT.scala 14:10]
  assign op_I_8_2_2 = I_8_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_9_1_2 = I_9_1_2; // @[MapT.scala 14:10]
  assign op_I_9_2_0 = I_9_2_0; // @[MapT.scala 14:10]
  assign op_I_9_2_1 = I_9_2_1; // @[MapT.scala 14:10]
  assign op_I_9_2_2 = I_9_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_10_1_2 = I_10_1_2; // @[MapT.scala 14:10]
  assign op_I_10_2_0 = I_10_2_0; // @[MapT.scala 14:10]
  assign op_I_10_2_1 = I_10_2_1; // @[MapT.scala 14:10]
  assign op_I_10_2_2 = I_10_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_11_1_2 = I_11_1_2; // @[MapT.scala 14:10]
  assign op_I_11_2_0 = I_11_2_0; // @[MapT.scala 14:10]
  assign op_I_11_2_1 = I_11_2_1; // @[MapT.scala 14:10]
  assign op_I_11_2_2 = I_11_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_12_1_2 = I_12_1_2; // @[MapT.scala 14:10]
  assign op_I_12_2_0 = I_12_2_0; // @[MapT.scala 14:10]
  assign op_I_12_2_1 = I_12_2_1; // @[MapT.scala 14:10]
  assign op_I_12_2_2 = I_12_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_13_1_2 = I_13_1_2; // @[MapT.scala 14:10]
  assign op_I_13_2_0 = I_13_2_0; // @[MapT.scala 14:10]
  assign op_I_13_2_1 = I_13_2_1; // @[MapT.scala 14:10]
  assign op_I_13_2_2 = I_13_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_14_1_2 = I_14_1_2; // @[MapT.scala 14:10]
  assign op_I_14_2_0 = I_14_2_0; // @[MapT.scala 14:10]
  assign op_I_14_2_1 = I_14_2_1; // @[MapT.scala 14:10]
  assign op_I_14_2_2 = I_14_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
  assign op_I_15_1_2 = I_15_1_2; // @[MapT.scala 14:10]
  assign op_I_15_2_0 = I_15_2_0; // @[MapT.scala 14:10]
  assign op_I_15_2_1 = I_15_2_1; // @[MapT.scala 14:10]
  assign op_I_15_2_2 = I_15_2_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [15:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_0_2,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_0_0_1_2,
  input  [15:0] I_0_0_2_0,
  input  [15:0] I_0_0_2_1,
  input  [15:0] I_0_0_2_2,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_0_2,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_1_0_1_2,
  input  [15:0] I_1_0_2_0,
  input  [15:0] I_1_0_2_1,
  input  [15:0] I_1_0_2_2,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_0_2,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_2_0_1_2,
  input  [15:0] I_2_0_2_0,
  input  [15:0] I_2_0_2_1,
  input  [15:0] I_2_0_2_2,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_0_2,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  input  [15:0] I_3_0_1_2,
  input  [15:0] I_3_0_2_0,
  input  [15:0] I_3_0_2_1,
  input  [15:0] I_3_0_2_2,
  input  [15:0] I_4_0_0_0,
  input  [15:0] I_4_0_0_1,
  input  [15:0] I_4_0_0_2,
  input  [15:0] I_4_0_1_0,
  input  [15:0] I_4_0_1_1,
  input  [15:0] I_4_0_1_2,
  input  [15:0] I_4_0_2_0,
  input  [15:0] I_4_0_2_1,
  input  [15:0] I_4_0_2_2,
  input  [15:0] I_5_0_0_0,
  input  [15:0] I_5_0_0_1,
  input  [15:0] I_5_0_0_2,
  input  [15:0] I_5_0_1_0,
  input  [15:0] I_5_0_1_1,
  input  [15:0] I_5_0_1_2,
  input  [15:0] I_5_0_2_0,
  input  [15:0] I_5_0_2_1,
  input  [15:0] I_5_0_2_2,
  input  [15:0] I_6_0_0_0,
  input  [15:0] I_6_0_0_1,
  input  [15:0] I_6_0_0_2,
  input  [15:0] I_6_0_1_0,
  input  [15:0] I_6_0_1_1,
  input  [15:0] I_6_0_1_2,
  input  [15:0] I_6_0_2_0,
  input  [15:0] I_6_0_2_1,
  input  [15:0] I_6_0_2_2,
  input  [15:0] I_7_0_0_0,
  input  [15:0] I_7_0_0_1,
  input  [15:0] I_7_0_0_2,
  input  [15:0] I_7_0_1_0,
  input  [15:0] I_7_0_1_1,
  input  [15:0] I_7_0_1_2,
  input  [15:0] I_7_0_2_0,
  input  [15:0] I_7_0_2_1,
  input  [15:0] I_7_0_2_2,
  input  [15:0] I_8_0_0_0,
  input  [15:0] I_8_0_0_1,
  input  [15:0] I_8_0_0_2,
  input  [15:0] I_8_0_1_0,
  input  [15:0] I_8_0_1_1,
  input  [15:0] I_8_0_1_2,
  input  [15:0] I_8_0_2_0,
  input  [15:0] I_8_0_2_1,
  input  [15:0] I_8_0_2_2,
  input  [15:0] I_9_0_0_0,
  input  [15:0] I_9_0_0_1,
  input  [15:0] I_9_0_0_2,
  input  [15:0] I_9_0_1_0,
  input  [15:0] I_9_0_1_1,
  input  [15:0] I_9_0_1_2,
  input  [15:0] I_9_0_2_0,
  input  [15:0] I_9_0_2_1,
  input  [15:0] I_9_0_2_2,
  input  [15:0] I_10_0_0_0,
  input  [15:0] I_10_0_0_1,
  input  [15:0] I_10_0_0_2,
  input  [15:0] I_10_0_1_0,
  input  [15:0] I_10_0_1_1,
  input  [15:0] I_10_0_1_2,
  input  [15:0] I_10_0_2_0,
  input  [15:0] I_10_0_2_1,
  input  [15:0] I_10_0_2_2,
  input  [15:0] I_11_0_0_0,
  input  [15:0] I_11_0_0_1,
  input  [15:0] I_11_0_0_2,
  input  [15:0] I_11_0_1_0,
  input  [15:0] I_11_0_1_1,
  input  [15:0] I_11_0_1_2,
  input  [15:0] I_11_0_2_0,
  input  [15:0] I_11_0_2_1,
  input  [15:0] I_11_0_2_2,
  input  [15:0] I_12_0_0_0,
  input  [15:0] I_12_0_0_1,
  input  [15:0] I_12_0_0_2,
  input  [15:0] I_12_0_1_0,
  input  [15:0] I_12_0_1_1,
  input  [15:0] I_12_0_1_2,
  input  [15:0] I_12_0_2_0,
  input  [15:0] I_12_0_2_1,
  input  [15:0] I_12_0_2_2,
  input  [15:0] I_13_0_0_0,
  input  [15:0] I_13_0_0_1,
  input  [15:0] I_13_0_0_2,
  input  [15:0] I_13_0_1_0,
  input  [15:0] I_13_0_1_1,
  input  [15:0] I_13_0_1_2,
  input  [15:0] I_13_0_2_0,
  input  [15:0] I_13_0_2_1,
  input  [15:0] I_13_0_2_2,
  input  [15:0] I_14_0_0_0,
  input  [15:0] I_14_0_0_1,
  input  [15:0] I_14_0_0_2,
  input  [15:0] I_14_0_1_0,
  input  [15:0] I_14_0_1_1,
  input  [15:0] I_14_0_1_2,
  input  [15:0] I_14_0_2_0,
  input  [15:0] I_14_0_2_1,
  input  [15:0] I_14_0_2_2,
  input  [15:0] I_15_0_0_0,
  input  [15:0] I_15_0_0_1,
  input  [15:0] I_15_0_0_2,
  input  [15:0] I_15_0_1_0,
  input  [15:0] I_15_0_1_1,
  input  [15:0] I_15_0_1_2,
  input  [15:0] I_15_0_2_0,
  input  [15:0] I_15_0_2_1,
  input  [15:0] I_15_0_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_8_1_0,
  output [15:0] O_8_1_1,
  output [15:0] O_8_1_2,
  output [15:0] O_8_2_0,
  output [15:0] O_8_2_1,
  output [15:0] O_8_2_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_9_1_0,
  output [15:0] O_9_1_1,
  output [15:0] O_9_1_2,
  output [15:0] O_9_2_0,
  output [15:0] O_9_2_1,
  output [15:0] O_9_2_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_10_1_0,
  output [15:0] O_10_1_1,
  output [15:0] O_10_1_2,
  output [15:0] O_10_2_0,
  output [15:0] O_10_2_1,
  output [15:0] O_10_2_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_11_1_0,
  output [15:0] O_11_1_1,
  output [15:0] O_11_1_2,
  output [15:0] O_11_2_0,
  output [15:0] O_11_2_1,
  output [15:0] O_11_2_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_12_1_0,
  output [15:0] O_12_1_1,
  output [15:0] O_12_1_2,
  output [15:0] O_12_2_0,
  output [15:0] O_12_2_1,
  output [15:0] O_12_2_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_13_1_0,
  output [15:0] O_13_1_1,
  output [15:0] O_13_1_2,
  output [15:0] O_13_2_0,
  output [15:0] O_13_2_1,
  output [15:0] O_13_2_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_14_1_0,
  output [15:0] O_14_1_1,
  output [15:0] O_14_1_2,
  output [15:0] O_14_2_0,
  output [15:0] O_14_2_1,
  output [15:0] O_14_2_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2,
  output [15:0] O_15_1_0,
  output [15:0] O_15_1_1,
  output [15:0] O_15_1_2,
  output [15:0] O_15_2_0,
  output [15:0] O_15_2_1,
  output [15:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  Remove1S_3 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0_0(other_ops_7_I_0_0_0),
    .I_0_0_1(other_ops_7_I_0_0_1),
    .I_0_0_2(other_ops_7_I_0_0_2),
    .I_0_1_0(other_ops_7_I_0_1_0),
    .I_0_1_1(other_ops_7_I_0_1_1),
    .I_0_1_2(other_ops_7_I_0_1_2),
    .I_0_2_0(other_ops_7_I_0_2_0),
    .I_0_2_1(other_ops_7_I_0_2_1),
    .I_0_2_2(other_ops_7_I_0_2_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  Remove1S_3 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0_0(other_ops_8_I_0_0_0),
    .I_0_0_1(other_ops_8_I_0_0_1),
    .I_0_0_2(other_ops_8_I_0_0_2),
    .I_0_1_0(other_ops_8_I_0_1_0),
    .I_0_1_1(other_ops_8_I_0_1_1),
    .I_0_1_2(other_ops_8_I_0_1_2),
    .I_0_2_0(other_ops_8_I_0_2_0),
    .I_0_2_1(other_ops_8_I_0_2_1),
    .I_0_2_2(other_ops_8_I_0_2_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  Remove1S_3 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0_0(other_ops_9_I_0_0_0),
    .I_0_0_1(other_ops_9_I_0_0_1),
    .I_0_0_2(other_ops_9_I_0_0_2),
    .I_0_1_0(other_ops_9_I_0_1_0),
    .I_0_1_1(other_ops_9_I_0_1_1),
    .I_0_1_2(other_ops_9_I_0_1_2),
    .I_0_2_0(other_ops_9_I_0_2_0),
    .I_0_2_1(other_ops_9_I_0_2_1),
    .I_0_2_2(other_ops_9_I_0_2_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  Remove1S_3 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0_0(other_ops_10_I_0_0_0),
    .I_0_0_1(other_ops_10_I_0_0_1),
    .I_0_0_2(other_ops_10_I_0_0_2),
    .I_0_1_0(other_ops_10_I_0_1_0),
    .I_0_1_1(other_ops_10_I_0_1_1),
    .I_0_1_2(other_ops_10_I_0_1_2),
    .I_0_2_0(other_ops_10_I_0_2_0),
    .I_0_2_1(other_ops_10_I_0_2_1),
    .I_0_2_2(other_ops_10_I_0_2_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  Remove1S_3 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0_0(other_ops_11_I_0_0_0),
    .I_0_0_1(other_ops_11_I_0_0_1),
    .I_0_0_2(other_ops_11_I_0_0_2),
    .I_0_1_0(other_ops_11_I_0_1_0),
    .I_0_1_1(other_ops_11_I_0_1_1),
    .I_0_1_2(other_ops_11_I_0_1_2),
    .I_0_2_0(other_ops_11_I_0_2_0),
    .I_0_2_1(other_ops_11_I_0_2_1),
    .I_0_2_2(other_ops_11_I_0_2_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  Remove1S_3 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0_0(other_ops_12_I_0_0_0),
    .I_0_0_1(other_ops_12_I_0_0_1),
    .I_0_0_2(other_ops_12_I_0_0_2),
    .I_0_1_0(other_ops_12_I_0_1_0),
    .I_0_1_1(other_ops_12_I_0_1_1),
    .I_0_1_2(other_ops_12_I_0_1_2),
    .I_0_2_0(other_ops_12_I_0_2_0),
    .I_0_2_1(other_ops_12_I_0_2_1),
    .I_0_2_2(other_ops_12_I_0_2_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  Remove1S_3 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0_0(other_ops_13_I_0_0_0),
    .I_0_0_1(other_ops_13_I_0_0_1),
    .I_0_0_2(other_ops_13_I_0_0_2),
    .I_0_1_0(other_ops_13_I_0_1_0),
    .I_0_1_1(other_ops_13_I_0_1_1),
    .I_0_1_2(other_ops_13_I_0_1_2),
    .I_0_2_0(other_ops_13_I_0_2_0),
    .I_0_2_1(other_ops_13_I_0_2_1),
    .I_0_2_2(other_ops_13_I_0_2_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  Remove1S_3 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0_0(other_ops_14_I_0_0_0),
    .I_0_0_1(other_ops_14_I_0_0_1),
    .I_0_0_2(other_ops_14_I_0_0_2),
    .I_0_1_0(other_ops_14_I_0_1_0),
    .I_0_1_1(other_ops_14_I_0_1_1),
    .I_0_1_2(other_ops_14_I_0_1_2),
    .I_0_2_0(other_ops_14_I_0_2_0),
    .I_0_2_1(other_ops_14_I_0_2_1),
    .I_0_2_2(other_ops_14_I_0_2_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[MapS.scala 21:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[MapS.scala 21:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[MapS.scala 21:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[MapS.scala 21:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[MapS.scala 21:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[MapS.scala 21:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[MapS.scala 21:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[MapS.scala 21:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[MapS.scala 21:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[MapS.scala 21:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[MapS.scala 21:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[MapS.scala 21:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[MapS.scala 21:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[MapS.scala 21:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[MapS.scala 21:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[MapS.scala 21:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[MapS.scala 21:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[MapS.scala 21:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[MapS.scala 21:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[MapS.scala 21:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[MapS.scala 21:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[MapS.scala 21:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[MapS.scala 21:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[MapS.scala 21:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[MapS.scala 21:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[MapS.scala 21:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[MapS.scala 21:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[MapS.scala 21:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[MapS.scala 21:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[MapS.scala 21:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[MapS.scala 21:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[MapS.scala 21:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[MapS.scala 21:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[MapS.scala 21:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[MapS.scala 21:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[MapS.scala 21:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[MapS.scala 21:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[MapS.scala 21:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[MapS.scala 21:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[MapS.scala 21:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[MapS.scala 21:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[MapS.scala 21:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[MapS.scala 21:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[MapS.scala 21:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[MapS.scala 21:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[MapS.scala 21:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[MapS.scala 21:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[MapS.scala 21:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[MapS.scala 21:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[MapS.scala 21:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[MapS.scala 21:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[MapS.scala 21:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[MapS.scala 21:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[MapS.scala 21:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[MapS.scala 21:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[MapS.scala 21:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0_0 = I_8_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_1 = I_8_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_2 = I_8_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_0 = I_8_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_1 = I_8_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_2 = I_8_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_0 = I_8_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_1 = I_8_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_2 = I_8_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0_0 = I_9_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_1 = I_9_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_2 = I_9_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_0 = I_9_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_1 = I_9_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_2 = I_9_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_0 = I_9_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_1 = I_9_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_2 = I_9_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0_0 = I_10_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_1 = I_10_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_2 = I_10_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_0 = I_10_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_1 = I_10_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_2 = I_10_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_0 = I_10_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_1 = I_10_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_2 = I_10_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0_0 = I_11_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_1 = I_11_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_2 = I_11_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_0 = I_11_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_1 = I_11_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_2 = I_11_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_0 = I_11_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_1 = I_11_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_2 = I_11_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0_0 = I_12_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_1 = I_12_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_2 = I_12_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_0 = I_12_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_1 = I_12_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_2 = I_12_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_0 = I_12_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_1 = I_12_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_2 = I_12_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0_0 = I_13_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_1 = I_13_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_2 = I_13_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_0 = I_13_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_1 = I_13_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_2 = I_13_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_0 = I_13_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_1 = I_13_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_2 = I_13_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0_0 = I_14_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_1 = I_14_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_2 = I_14_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_0 = I_14_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_1 = I_14_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_2 = I_14_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_0 = I_14_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_1 = I_14_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_2 = I_14_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0_0 = I_15_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_1 = I_15_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_2 = I_15_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_0 = I_15_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_1 = I_15_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_2 = I_15_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_0 = I_15_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_1 = I_15_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_2 = I_15_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0_0,
  input  [15:0] I_0_0_0_1,
  input  [15:0] I_0_0_0_2,
  input  [15:0] I_0_0_1_0,
  input  [15:0] I_0_0_1_1,
  input  [15:0] I_0_0_1_2,
  input  [15:0] I_0_0_2_0,
  input  [15:0] I_0_0_2_1,
  input  [15:0] I_0_0_2_2,
  input  [15:0] I_1_0_0_0,
  input  [15:0] I_1_0_0_1,
  input  [15:0] I_1_0_0_2,
  input  [15:0] I_1_0_1_0,
  input  [15:0] I_1_0_1_1,
  input  [15:0] I_1_0_1_2,
  input  [15:0] I_1_0_2_0,
  input  [15:0] I_1_0_2_1,
  input  [15:0] I_1_0_2_2,
  input  [15:0] I_2_0_0_0,
  input  [15:0] I_2_0_0_1,
  input  [15:0] I_2_0_0_2,
  input  [15:0] I_2_0_1_0,
  input  [15:0] I_2_0_1_1,
  input  [15:0] I_2_0_1_2,
  input  [15:0] I_2_0_2_0,
  input  [15:0] I_2_0_2_1,
  input  [15:0] I_2_0_2_2,
  input  [15:0] I_3_0_0_0,
  input  [15:0] I_3_0_0_1,
  input  [15:0] I_3_0_0_2,
  input  [15:0] I_3_0_1_0,
  input  [15:0] I_3_0_1_1,
  input  [15:0] I_3_0_1_2,
  input  [15:0] I_3_0_2_0,
  input  [15:0] I_3_0_2_1,
  input  [15:0] I_3_0_2_2,
  input  [15:0] I_4_0_0_0,
  input  [15:0] I_4_0_0_1,
  input  [15:0] I_4_0_0_2,
  input  [15:0] I_4_0_1_0,
  input  [15:0] I_4_0_1_1,
  input  [15:0] I_4_0_1_2,
  input  [15:0] I_4_0_2_0,
  input  [15:0] I_4_0_2_1,
  input  [15:0] I_4_0_2_2,
  input  [15:0] I_5_0_0_0,
  input  [15:0] I_5_0_0_1,
  input  [15:0] I_5_0_0_2,
  input  [15:0] I_5_0_1_0,
  input  [15:0] I_5_0_1_1,
  input  [15:0] I_5_0_1_2,
  input  [15:0] I_5_0_2_0,
  input  [15:0] I_5_0_2_1,
  input  [15:0] I_5_0_2_2,
  input  [15:0] I_6_0_0_0,
  input  [15:0] I_6_0_0_1,
  input  [15:0] I_6_0_0_2,
  input  [15:0] I_6_0_1_0,
  input  [15:0] I_6_0_1_1,
  input  [15:0] I_6_0_1_2,
  input  [15:0] I_6_0_2_0,
  input  [15:0] I_6_0_2_1,
  input  [15:0] I_6_0_2_2,
  input  [15:0] I_7_0_0_0,
  input  [15:0] I_7_0_0_1,
  input  [15:0] I_7_0_0_2,
  input  [15:0] I_7_0_1_0,
  input  [15:0] I_7_0_1_1,
  input  [15:0] I_7_0_1_2,
  input  [15:0] I_7_0_2_0,
  input  [15:0] I_7_0_2_1,
  input  [15:0] I_7_0_2_2,
  input  [15:0] I_8_0_0_0,
  input  [15:0] I_8_0_0_1,
  input  [15:0] I_8_0_0_2,
  input  [15:0] I_8_0_1_0,
  input  [15:0] I_8_0_1_1,
  input  [15:0] I_8_0_1_2,
  input  [15:0] I_8_0_2_0,
  input  [15:0] I_8_0_2_1,
  input  [15:0] I_8_0_2_2,
  input  [15:0] I_9_0_0_0,
  input  [15:0] I_9_0_0_1,
  input  [15:0] I_9_0_0_2,
  input  [15:0] I_9_0_1_0,
  input  [15:0] I_9_0_1_1,
  input  [15:0] I_9_0_1_2,
  input  [15:0] I_9_0_2_0,
  input  [15:0] I_9_0_2_1,
  input  [15:0] I_9_0_2_2,
  input  [15:0] I_10_0_0_0,
  input  [15:0] I_10_0_0_1,
  input  [15:0] I_10_0_0_2,
  input  [15:0] I_10_0_1_0,
  input  [15:0] I_10_0_1_1,
  input  [15:0] I_10_0_1_2,
  input  [15:0] I_10_0_2_0,
  input  [15:0] I_10_0_2_1,
  input  [15:0] I_10_0_2_2,
  input  [15:0] I_11_0_0_0,
  input  [15:0] I_11_0_0_1,
  input  [15:0] I_11_0_0_2,
  input  [15:0] I_11_0_1_0,
  input  [15:0] I_11_0_1_1,
  input  [15:0] I_11_0_1_2,
  input  [15:0] I_11_0_2_0,
  input  [15:0] I_11_0_2_1,
  input  [15:0] I_11_0_2_2,
  input  [15:0] I_12_0_0_0,
  input  [15:0] I_12_0_0_1,
  input  [15:0] I_12_0_0_2,
  input  [15:0] I_12_0_1_0,
  input  [15:0] I_12_0_1_1,
  input  [15:0] I_12_0_1_2,
  input  [15:0] I_12_0_2_0,
  input  [15:0] I_12_0_2_1,
  input  [15:0] I_12_0_2_2,
  input  [15:0] I_13_0_0_0,
  input  [15:0] I_13_0_0_1,
  input  [15:0] I_13_0_0_2,
  input  [15:0] I_13_0_1_0,
  input  [15:0] I_13_0_1_1,
  input  [15:0] I_13_0_1_2,
  input  [15:0] I_13_0_2_0,
  input  [15:0] I_13_0_2_1,
  input  [15:0] I_13_0_2_2,
  input  [15:0] I_14_0_0_0,
  input  [15:0] I_14_0_0_1,
  input  [15:0] I_14_0_0_2,
  input  [15:0] I_14_0_1_0,
  input  [15:0] I_14_0_1_1,
  input  [15:0] I_14_0_1_2,
  input  [15:0] I_14_0_2_0,
  input  [15:0] I_14_0_2_1,
  input  [15:0] I_14_0_2_2,
  input  [15:0] I_15_0_0_0,
  input  [15:0] I_15_0_0_1,
  input  [15:0] I_15_0_0_2,
  input  [15:0] I_15_0_1_0,
  input  [15:0] I_15_0_1_1,
  input  [15:0] I_15_0_1_2,
  input  [15:0] I_15_0_2_0,
  input  [15:0] I_15_0_2_1,
  input  [15:0] I_15_0_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_0_0_1,
  output [15:0] O_0_0_2,
  output [15:0] O_0_1_0,
  output [15:0] O_0_1_1,
  output [15:0] O_0_1_2,
  output [15:0] O_0_2_0,
  output [15:0] O_0_2_1,
  output [15:0] O_0_2_2,
  output [15:0] O_1_0_0,
  output [15:0] O_1_0_1,
  output [15:0] O_1_0_2,
  output [15:0] O_1_1_0,
  output [15:0] O_1_1_1,
  output [15:0] O_1_1_2,
  output [15:0] O_1_2_0,
  output [15:0] O_1_2_1,
  output [15:0] O_1_2_2,
  output [15:0] O_2_0_0,
  output [15:0] O_2_0_1,
  output [15:0] O_2_0_2,
  output [15:0] O_2_1_0,
  output [15:0] O_2_1_1,
  output [15:0] O_2_1_2,
  output [15:0] O_2_2_0,
  output [15:0] O_2_2_1,
  output [15:0] O_2_2_2,
  output [15:0] O_3_0_0,
  output [15:0] O_3_0_1,
  output [15:0] O_3_0_2,
  output [15:0] O_3_1_0,
  output [15:0] O_3_1_1,
  output [15:0] O_3_1_2,
  output [15:0] O_3_2_0,
  output [15:0] O_3_2_1,
  output [15:0] O_3_2_2,
  output [15:0] O_4_0_0,
  output [15:0] O_4_0_1,
  output [15:0] O_4_0_2,
  output [15:0] O_4_1_0,
  output [15:0] O_4_1_1,
  output [15:0] O_4_1_2,
  output [15:0] O_4_2_0,
  output [15:0] O_4_2_1,
  output [15:0] O_4_2_2,
  output [15:0] O_5_0_0,
  output [15:0] O_5_0_1,
  output [15:0] O_5_0_2,
  output [15:0] O_5_1_0,
  output [15:0] O_5_1_1,
  output [15:0] O_5_1_2,
  output [15:0] O_5_2_0,
  output [15:0] O_5_2_1,
  output [15:0] O_5_2_2,
  output [15:0] O_6_0_0,
  output [15:0] O_6_0_1,
  output [15:0] O_6_0_2,
  output [15:0] O_6_1_0,
  output [15:0] O_6_1_1,
  output [15:0] O_6_1_2,
  output [15:0] O_6_2_0,
  output [15:0] O_6_2_1,
  output [15:0] O_6_2_2,
  output [15:0] O_7_0_0,
  output [15:0] O_7_0_1,
  output [15:0] O_7_0_2,
  output [15:0] O_7_1_0,
  output [15:0] O_7_1_1,
  output [15:0] O_7_1_2,
  output [15:0] O_7_2_0,
  output [15:0] O_7_2_1,
  output [15:0] O_7_2_2,
  output [15:0] O_8_0_0,
  output [15:0] O_8_0_1,
  output [15:0] O_8_0_2,
  output [15:0] O_8_1_0,
  output [15:0] O_8_1_1,
  output [15:0] O_8_1_2,
  output [15:0] O_8_2_0,
  output [15:0] O_8_2_1,
  output [15:0] O_8_2_2,
  output [15:0] O_9_0_0,
  output [15:0] O_9_0_1,
  output [15:0] O_9_0_2,
  output [15:0] O_9_1_0,
  output [15:0] O_9_1_1,
  output [15:0] O_9_1_2,
  output [15:0] O_9_2_0,
  output [15:0] O_9_2_1,
  output [15:0] O_9_2_2,
  output [15:0] O_10_0_0,
  output [15:0] O_10_0_1,
  output [15:0] O_10_0_2,
  output [15:0] O_10_1_0,
  output [15:0] O_10_1_1,
  output [15:0] O_10_1_2,
  output [15:0] O_10_2_0,
  output [15:0] O_10_2_1,
  output [15:0] O_10_2_2,
  output [15:0] O_11_0_0,
  output [15:0] O_11_0_1,
  output [15:0] O_11_0_2,
  output [15:0] O_11_1_0,
  output [15:0] O_11_1_1,
  output [15:0] O_11_1_2,
  output [15:0] O_11_2_0,
  output [15:0] O_11_2_1,
  output [15:0] O_11_2_2,
  output [15:0] O_12_0_0,
  output [15:0] O_12_0_1,
  output [15:0] O_12_0_2,
  output [15:0] O_12_1_0,
  output [15:0] O_12_1_1,
  output [15:0] O_12_1_2,
  output [15:0] O_12_2_0,
  output [15:0] O_12_2_1,
  output [15:0] O_12_2_2,
  output [15:0] O_13_0_0,
  output [15:0] O_13_0_1,
  output [15:0] O_13_0_2,
  output [15:0] O_13_1_0,
  output [15:0] O_13_1_1,
  output [15:0] O_13_1_2,
  output [15:0] O_13_2_0,
  output [15:0] O_13_2_1,
  output [15:0] O_13_2_2,
  output [15:0] O_14_0_0,
  output [15:0] O_14_0_1,
  output [15:0] O_14_0_2,
  output [15:0] O_14_1_0,
  output [15:0] O_14_1_1,
  output [15:0] O_14_1_2,
  output [15:0] O_14_2_0,
  output [15:0] O_14_2_1,
  output [15:0] O_14_2_2,
  output [15:0] O_15_0_0,
  output [15:0] O_15_0_1,
  output [15:0] O_15_0_2,
  output [15:0] O_15_1_0,
  output [15:0] O_15_1_1,
  output [15:0] O_15_1_2,
  output [15:0] O_15_2_0,
  output [15:0] O_15_2_1,
  output [15:0] O_15_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_2_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_4_0_1_2(op_I_4_0_1_2),
    .I_4_0_2_0(op_I_4_0_2_0),
    .I_4_0_2_1(op_I_4_0_2_1),
    .I_4_0_2_2(op_I_4_0_2_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_5_0_1_2(op_I_5_0_1_2),
    .I_5_0_2_0(op_I_5_0_2_0),
    .I_5_0_2_1(op_I_5_0_2_1),
    .I_5_0_2_2(op_I_5_0_2_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_6_0_1_2(op_I_6_0_1_2),
    .I_6_0_2_0(op_I_6_0_2_0),
    .I_6_0_2_1(op_I_6_0_2_1),
    .I_6_0_2_2(op_I_6_0_2_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_7_0_1_2(op_I_7_0_1_2),
    .I_7_0_2_0(op_I_7_0_2_0),
    .I_7_0_2_1(op_I_7_0_2_1),
    .I_7_0_2_2(op_I_7_0_2_2),
    .I_8_0_0_0(op_I_8_0_0_0),
    .I_8_0_0_1(op_I_8_0_0_1),
    .I_8_0_0_2(op_I_8_0_0_2),
    .I_8_0_1_0(op_I_8_0_1_0),
    .I_8_0_1_1(op_I_8_0_1_1),
    .I_8_0_1_2(op_I_8_0_1_2),
    .I_8_0_2_0(op_I_8_0_2_0),
    .I_8_0_2_1(op_I_8_0_2_1),
    .I_8_0_2_2(op_I_8_0_2_2),
    .I_9_0_0_0(op_I_9_0_0_0),
    .I_9_0_0_1(op_I_9_0_0_1),
    .I_9_0_0_2(op_I_9_0_0_2),
    .I_9_0_1_0(op_I_9_0_1_0),
    .I_9_0_1_1(op_I_9_0_1_1),
    .I_9_0_1_2(op_I_9_0_1_2),
    .I_9_0_2_0(op_I_9_0_2_0),
    .I_9_0_2_1(op_I_9_0_2_1),
    .I_9_0_2_2(op_I_9_0_2_2),
    .I_10_0_0_0(op_I_10_0_0_0),
    .I_10_0_0_1(op_I_10_0_0_1),
    .I_10_0_0_2(op_I_10_0_0_2),
    .I_10_0_1_0(op_I_10_0_1_0),
    .I_10_0_1_1(op_I_10_0_1_1),
    .I_10_0_1_2(op_I_10_0_1_2),
    .I_10_0_2_0(op_I_10_0_2_0),
    .I_10_0_2_1(op_I_10_0_2_1),
    .I_10_0_2_2(op_I_10_0_2_2),
    .I_11_0_0_0(op_I_11_0_0_0),
    .I_11_0_0_1(op_I_11_0_0_1),
    .I_11_0_0_2(op_I_11_0_0_2),
    .I_11_0_1_0(op_I_11_0_1_0),
    .I_11_0_1_1(op_I_11_0_1_1),
    .I_11_0_1_2(op_I_11_0_1_2),
    .I_11_0_2_0(op_I_11_0_2_0),
    .I_11_0_2_1(op_I_11_0_2_1),
    .I_11_0_2_2(op_I_11_0_2_2),
    .I_12_0_0_0(op_I_12_0_0_0),
    .I_12_0_0_1(op_I_12_0_0_1),
    .I_12_0_0_2(op_I_12_0_0_2),
    .I_12_0_1_0(op_I_12_0_1_0),
    .I_12_0_1_1(op_I_12_0_1_1),
    .I_12_0_1_2(op_I_12_0_1_2),
    .I_12_0_2_0(op_I_12_0_2_0),
    .I_12_0_2_1(op_I_12_0_2_1),
    .I_12_0_2_2(op_I_12_0_2_2),
    .I_13_0_0_0(op_I_13_0_0_0),
    .I_13_0_0_1(op_I_13_0_0_1),
    .I_13_0_0_2(op_I_13_0_0_2),
    .I_13_0_1_0(op_I_13_0_1_0),
    .I_13_0_1_1(op_I_13_0_1_1),
    .I_13_0_1_2(op_I_13_0_1_2),
    .I_13_0_2_0(op_I_13_0_2_0),
    .I_13_0_2_1(op_I_13_0_2_1),
    .I_13_0_2_2(op_I_13_0_2_2),
    .I_14_0_0_0(op_I_14_0_0_0),
    .I_14_0_0_1(op_I_14_0_0_1),
    .I_14_0_0_2(op_I_14_0_0_2),
    .I_14_0_1_0(op_I_14_0_1_0),
    .I_14_0_1_1(op_I_14_0_1_1),
    .I_14_0_1_2(op_I_14_0_1_2),
    .I_14_0_2_0(op_I_14_0_2_0),
    .I_14_0_2_1(op_I_14_0_2_1),
    .I_14_0_2_2(op_I_14_0_2_2),
    .I_15_0_0_0(op_I_15_0_0_0),
    .I_15_0_0_1(op_I_15_0_0_1),
    .I_15_0_0_2(op_I_15_0_0_2),
    .I_15_0_1_0(op_I_15_0_1_0),
    .I_15_0_1_1(op_I_15_0_1_1),
    .I_15_0_1_2(op_I_15_0_1_2),
    .I_15_0_2_0(op_I_15_0_2_0),
    .I_15_0_2_1(op_I_15_0_2_1),
    .I_15_0_2_2(op_I_15_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_8_2_0(op_O_8_2_0),
    .O_8_2_1(op_O_8_2_1),
    .O_8_2_2(op_O_8_2_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_9_2_0(op_O_9_2_0),
    .O_9_2_1(op_O_9_2_1),
    .O_9_2_2(op_O_9_2_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_10_2_0(op_O_10_2_0),
    .O_10_2_1(op_O_10_2_1),
    .O_10_2_2(op_O_10_2_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_11_2_0(op_O_11_2_0),
    .O_11_2_1(op_O_11_2_1),
    .O_11_2_2(op_O_11_2_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_12_2_0(op_O_12_2_0),
    .O_12_2_1(op_O_12_2_1),
    .O_12_2_2(op_O_12_2_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_13_2_0(op_O_13_2_0),
    .O_13_2_1(op_O_13_2_1),
    .O_13_2_2(op_O_13_2_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_14_2_0(op_O_14_2_0),
    .O_14_2_1(op_O_14_2_1),
    .O_14_2_2(op_O_14_2_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2),
    .O_15_2_0(op_O_15_2_0),
    .O_15_2_1(op_O_15_2_1),
    .O_15_2_2(op_O_15_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_4_1_2 = op_O_4_1_2; // @[MapT.scala 15:7]
  assign O_4_2_0 = op_O_4_2_0; // @[MapT.scala 15:7]
  assign O_4_2_1 = op_O_4_2_1; // @[MapT.scala 15:7]
  assign O_4_2_2 = op_O_4_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_5_1_2 = op_O_5_1_2; // @[MapT.scala 15:7]
  assign O_5_2_0 = op_O_5_2_0; // @[MapT.scala 15:7]
  assign O_5_2_1 = op_O_5_2_1; // @[MapT.scala 15:7]
  assign O_5_2_2 = op_O_5_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_6_1_2 = op_O_6_1_2; // @[MapT.scala 15:7]
  assign O_6_2_0 = op_O_6_2_0; // @[MapT.scala 15:7]
  assign O_6_2_1 = op_O_6_2_1; // @[MapT.scala 15:7]
  assign O_6_2_2 = op_O_6_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_7_1_2 = op_O_7_1_2; // @[MapT.scala 15:7]
  assign O_7_2_0 = op_O_7_2_0; // @[MapT.scala 15:7]
  assign O_7_2_1 = op_O_7_2_1; // @[MapT.scala 15:7]
  assign O_7_2_2 = op_O_7_2_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_8_1_0 = op_O_8_1_0; // @[MapT.scala 15:7]
  assign O_8_1_1 = op_O_8_1_1; // @[MapT.scala 15:7]
  assign O_8_1_2 = op_O_8_1_2; // @[MapT.scala 15:7]
  assign O_8_2_0 = op_O_8_2_0; // @[MapT.scala 15:7]
  assign O_8_2_1 = op_O_8_2_1; // @[MapT.scala 15:7]
  assign O_8_2_2 = op_O_8_2_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_9_1_0 = op_O_9_1_0; // @[MapT.scala 15:7]
  assign O_9_1_1 = op_O_9_1_1; // @[MapT.scala 15:7]
  assign O_9_1_2 = op_O_9_1_2; // @[MapT.scala 15:7]
  assign O_9_2_0 = op_O_9_2_0; // @[MapT.scala 15:7]
  assign O_9_2_1 = op_O_9_2_1; // @[MapT.scala 15:7]
  assign O_9_2_2 = op_O_9_2_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_10_1_0 = op_O_10_1_0; // @[MapT.scala 15:7]
  assign O_10_1_1 = op_O_10_1_1; // @[MapT.scala 15:7]
  assign O_10_1_2 = op_O_10_1_2; // @[MapT.scala 15:7]
  assign O_10_2_0 = op_O_10_2_0; // @[MapT.scala 15:7]
  assign O_10_2_1 = op_O_10_2_1; // @[MapT.scala 15:7]
  assign O_10_2_2 = op_O_10_2_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_11_1_0 = op_O_11_1_0; // @[MapT.scala 15:7]
  assign O_11_1_1 = op_O_11_1_1; // @[MapT.scala 15:7]
  assign O_11_1_2 = op_O_11_1_2; // @[MapT.scala 15:7]
  assign O_11_2_0 = op_O_11_2_0; // @[MapT.scala 15:7]
  assign O_11_2_1 = op_O_11_2_1; // @[MapT.scala 15:7]
  assign O_11_2_2 = op_O_11_2_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_12_1_0 = op_O_12_1_0; // @[MapT.scala 15:7]
  assign O_12_1_1 = op_O_12_1_1; // @[MapT.scala 15:7]
  assign O_12_1_2 = op_O_12_1_2; // @[MapT.scala 15:7]
  assign O_12_2_0 = op_O_12_2_0; // @[MapT.scala 15:7]
  assign O_12_2_1 = op_O_12_2_1; // @[MapT.scala 15:7]
  assign O_12_2_2 = op_O_12_2_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_13_1_0 = op_O_13_1_0; // @[MapT.scala 15:7]
  assign O_13_1_1 = op_O_13_1_1; // @[MapT.scala 15:7]
  assign O_13_1_2 = op_O_13_1_2; // @[MapT.scala 15:7]
  assign O_13_2_0 = op_O_13_2_0; // @[MapT.scala 15:7]
  assign O_13_2_1 = op_O_13_2_1; // @[MapT.scala 15:7]
  assign O_13_2_2 = op_O_13_2_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_14_1_0 = op_O_14_1_0; // @[MapT.scala 15:7]
  assign O_14_1_1 = op_O_14_1_1; // @[MapT.scala 15:7]
  assign O_14_1_2 = op_O_14_1_2; // @[MapT.scala 15:7]
  assign O_14_2_0 = op_O_14_2_0; // @[MapT.scala 15:7]
  assign O_14_2_1 = op_O_14_2_1; // @[MapT.scala 15:7]
  assign O_14_2_2 = op_O_14_2_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign O_15_1_0 = op_O_15_1_0; // @[MapT.scala 15:7]
  assign O_15_1_1 = op_O_15_1_1; // @[MapT.scala 15:7]
  assign O_15_1_2 = op_O_15_1_2; // @[MapT.scala 15:7]
  assign O_15_2_0 = op_O_15_2_0; // @[MapT.scala 15:7]
  assign O_15_2_1 = op_O_15_2_1; // @[MapT.scala 15:7]
  assign O_15_2_2 = op_O_15_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_2 = I_4_0_1_2; // @[MapT.scala 14:10]
  assign op_I_4_0_2_0 = I_4_0_2_0; // @[MapT.scala 14:10]
  assign op_I_4_0_2_1 = I_4_0_2_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2_2 = I_4_0_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_2 = I_5_0_1_2; // @[MapT.scala 14:10]
  assign op_I_5_0_2_0 = I_5_0_2_0; // @[MapT.scala 14:10]
  assign op_I_5_0_2_1 = I_5_0_2_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2_2 = I_5_0_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_2 = I_6_0_1_2; // @[MapT.scala 14:10]
  assign op_I_6_0_2_0 = I_6_0_2_0; // @[MapT.scala 14:10]
  assign op_I_6_0_2_1 = I_6_0_2_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2_2 = I_6_0_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_2 = I_7_0_1_2; // @[MapT.scala 14:10]
  assign op_I_7_0_2_0 = I_7_0_2_0; // @[MapT.scala 14:10]
  assign op_I_7_0_2_1 = I_7_0_2_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2_2 = I_7_0_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0_0 = I_8_0_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_0_1 = I_8_0_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0_2 = I_8_0_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_1_0 = I_8_0_1_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1_1 = I_8_0_1_1; // @[MapT.scala 14:10]
  assign op_I_8_0_1_2 = I_8_0_1_2; // @[MapT.scala 14:10]
  assign op_I_8_0_2_0 = I_8_0_2_0; // @[MapT.scala 14:10]
  assign op_I_8_0_2_1 = I_8_0_2_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2_2 = I_8_0_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0_0 = I_9_0_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_0_1 = I_9_0_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0_2 = I_9_0_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_1_0 = I_9_0_1_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1_1 = I_9_0_1_1; // @[MapT.scala 14:10]
  assign op_I_9_0_1_2 = I_9_0_1_2; // @[MapT.scala 14:10]
  assign op_I_9_0_2_0 = I_9_0_2_0; // @[MapT.scala 14:10]
  assign op_I_9_0_2_1 = I_9_0_2_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2_2 = I_9_0_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0_0 = I_10_0_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_0_1 = I_10_0_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0_2 = I_10_0_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_1_0 = I_10_0_1_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1_1 = I_10_0_1_1; // @[MapT.scala 14:10]
  assign op_I_10_0_1_2 = I_10_0_1_2; // @[MapT.scala 14:10]
  assign op_I_10_0_2_0 = I_10_0_2_0; // @[MapT.scala 14:10]
  assign op_I_10_0_2_1 = I_10_0_2_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2_2 = I_10_0_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0_0 = I_11_0_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_0_1 = I_11_0_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0_2 = I_11_0_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_1_0 = I_11_0_1_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1_1 = I_11_0_1_1; // @[MapT.scala 14:10]
  assign op_I_11_0_1_2 = I_11_0_1_2; // @[MapT.scala 14:10]
  assign op_I_11_0_2_0 = I_11_0_2_0; // @[MapT.scala 14:10]
  assign op_I_11_0_2_1 = I_11_0_2_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2_2 = I_11_0_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0_0 = I_12_0_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_0_1 = I_12_0_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0_2 = I_12_0_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_1_0 = I_12_0_1_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1_1 = I_12_0_1_1; // @[MapT.scala 14:10]
  assign op_I_12_0_1_2 = I_12_0_1_2; // @[MapT.scala 14:10]
  assign op_I_12_0_2_0 = I_12_0_2_0; // @[MapT.scala 14:10]
  assign op_I_12_0_2_1 = I_12_0_2_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2_2 = I_12_0_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0_0 = I_13_0_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_0_1 = I_13_0_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0_2 = I_13_0_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_1_0 = I_13_0_1_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1_1 = I_13_0_1_1; // @[MapT.scala 14:10]
  assign op_I_13_0_1_2 = I_13_0_1_2; // @[MapT.scala 14:10]
  assign op_I_13_0_2_0 = I_13_0_2_0; // @[MapT.scala 14:10]
  assign op_I_13_0_2_1 = I_13_0_2_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2_2 = I_13_0_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0_0 = I_14_0_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_0_1 = I_14_0_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0_2 = I_14_0_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_1_0 = I_14_0_1_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1_1 = I_14_0_1_1; // @[MapT.scala 14:10]
  assign op_I_14_0_1_2 = I_14_0_1_2; // @[MapT.scala 14:10]
  assign op_I_14_0_2_0 = I_14_0_2_0; // @[MapT.scala 14:10]
  assign op_I_14_0_2_1 = I_14_0_2_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2_2 = I_14_0_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0_0 = I_15_0_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_0_1 = I_15_0_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0_2 = I_15_0_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_1_0 = I_15_0_1_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1_1 = I_15_0_1_1; // @[MapT.scala 14:10]
  assign op_I_15_0_1_2 = I_15_0_1_2; // @[MapT.scala 14:10]
  assign op_I_15_0_2_0 = I_15_0_2_0; // @[MapT.scala 14:10]
  assign op_I_15_0_2_1 = I_15_0_2_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2_2 = I_15_0_2_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [2:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [2:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 3'h5; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 3'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 3'h5; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0,
  input  [7:0]  I1,
  output [15:0] O_t0b,
  output [7:0]  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  input  [15:0] I0_1,
  input  [15:0] I0_2,
  input  [7:0]  I1_0,
  input  [7:0]  I1_1,
  input  [7:0]  I1_2,
  output [15:0] O_0_t0b,
  output [7:0]  O_0_t1b,
  output [15:0] O_1_t0b,
  output [7:0]  O_1_t1b,
  output [15:0] O_2_t0b,
  output [7:0]  O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_9(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  input  [15:0] I0_0_1,
  input  [15:0] I0_0_2,
  input  [15:0] I0_1_0,
  input  [15:0] I0_1_1,
  input  [15:0] I0_1_2,
  input  [15:0] I0_2_0,
  input  [15:0] I0_2_1,
  input  [15:0] I0_2_2,
  output [15:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b,
  output [15:0] O_0_1_t0b,
  output [7:0]  O_0_1_t1b,
  output [15:0] O_0_2_t0b,
  output [7:0]  O_0_2_t1b,
  output [15:0] O_1_0_t0b,
  output [7:0]  O_1_0_t1b,
  output [15:0] O_1_1_t0b,
  output [7:0]  O_1_1_t1b,
  output [15:0] O_1_2_t0b,
  output [7:0]  O_1_2_t1b,
  output [15:0] O_2_0_t0b,
  output [7:0]  O_2_0_t1b,
  output [15:0] O_2_1_t0b,
  output [7:0]  O_2_1_t1b,
  output [15:0] O_2_2_t0b,
  output [7:0]  O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [15:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_8 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_8 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_8 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 8'h0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 8'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 8'h0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 8'h0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 8'h0; // @[Map2S.scala 23:43]
endmodule
module LShift(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_t0b,
  input  [7:0]  I_t1b,
  output [15:0] O
);
  wire [270:0] _GEN_0; // @[Arithmetic.scala 431:25]
  wire [270:0] _T; // @[Arithmetic.scala 431:25]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 431:25]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 431:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 433:14]
  assign O = _T[15:0]; // @[Arithmetic.scala 431:7]
endmodule
module MapS_4(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_t0b,
  input  [7:0]  I_0_t1b,
  input  [15:0] I_1_t0b,
  input  [7:0]  I_1_t1b,
  input  [15:0] I_2_t0b,
  input  [7:0]  I_2_t1b,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  LShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  LShift other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  LShift other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_5(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_t0b,
  input  [7:0]  I_0_0_t1b,
  input  [15:0] I_0_1_t0b,
  input  [7:0]  I_0_1_t1b,
  input  [15:0] I_0_2_t0b,
  input  [7:0]  I_0_2_t1b,
  input  [15:0] I_1_0_t0b,
  input  [7:0]  I_1_0_t1b,
  input  [15:0] I_1_1_t0b,
  input  [7:0]  I_1_1_t1b,
  input  [15:0] I_1_2_t0b,
  input  [7:0]  I_1_2_t1b,
  input  [15:0] I_2_0_t0b,
  input  [7:0]  I_2_0_t1b,
  input  [15:0] I_2_1_t0b,
  input  [7:0]  I_2_1_t1b,
  input  [15:0] I_2_2_t0b,
  input  [7:0]  I_2_2_t1b,
  output [15:0] O_0_0,
  output [15:0] O_0_1,
  output [15:0] O_0_2,
  output [15:0] O_1_0,
  output [15:0] O_1_1,
  output [15:0] O_1_2,
  output [15:0] O_2_0,
  output [15:0] O_2_1,
  output [15:0] O_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_4 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_4 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [15:0] I_t0b,
  input  [15:0] I_t1b,
  output [15:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  output [15:0] O_0
);
  wire [15:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [15:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = I_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = I_0; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = I_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module MapS_6(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0,
  output [15:0] O_1_0,
  output [15:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [15:0] I_0_t0b,
  input  [15:0] I_0_t1b,
  output [15:0] O_0
);
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [15:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [15:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_1_0,
  input  [15:0] I_2_0,
  output [15:0] O_0_0
);
  wire [15:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [15:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [15:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = I_0_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = I_1_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = I_2_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [2:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [2:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 3'h7; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 3'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 3'h7; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2S_10(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0,
  output [15:0] O_0_t0b,
  output [7:0]  O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = 8'h4; // @[Map2S.scala 18:13]
endmodule
module Map2S_11(
  input         valid_up,
  output        valid_down,
  input  [15:0] I0_0_0,
  output [15:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [15:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
endmodule
module RShift(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_t0b,
  input  [7:0]  I_t1b,
  output [15:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 402:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 400:7]
endmodule
module MapS_7(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_t0b,
  input  [7:0]  I_0_t1b,
  output [15:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O; // @[MapS.scala 9:22]
  RShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_8(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_t0b,
  input  [7:0]  I_0_0_t1b,
  output [15:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_0_1,
  input  [15:0] I_0_2,
  input  [15:0] I_1_0,
  input  [15:0] I_1_1,
  input  [15:0] I_1_2,
  input  [15:0] I_2_0,
  input  [15:0] I_2_1,
  input  [15:0] I_2_2,
  output [15:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n118_valid_up; // @[Top.scala 18:22]
  wire  n118_valid_down; // @[Top.scala 18:22]
  wire [15:0] n118_I0_0_0; // @[Top.scala 18:22]
  wire [15:0] n118_I0_0_1; // @[Top.scala 18:22]
  wire [15:0] n118_I0_0_2; // @[Top.scala 18:22]
  wire [15:0] n118_I0_1_0; // @[Top.scala 18:22]
  wire [15:0] n118_I0_1_1; // @[Top.scala 18:22]
  wire [15:0] n118_I0_1_2; // @[Top.scala 18:22]
  wire [15:0] n118_I0_2_0; // @[Top.scala 18:22]
  wire [15:0] n118_I0_2_1; // @[Top.scala 18:22]
  wire [15:0] n118_I0_2_2; // @[Top.scala 18:22]
  wire [15:0] n118_O_0_0_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_0_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_0_1_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_0_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_0_2_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_0_2_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_1_0_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_1_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_1_1_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_1_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_1_2_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_1_2_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_2_0_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_2_0_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_2_1_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_2_1_t1b; // @[Top.scala 18:22]
  wire [15:0] n118_O_2_2_t0b; // @[Top.scala 18:22]
  wire [7:0] n118_O_2_2_t1b; // @[Top.scala 18:22]
  wire  n129_valid_up; // @[Top.scala 22:22]
  wire  n129_valid_down; // @[Top.scala 22:22]
  wire [15:0] n129_I_0_0_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_0_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_0_1_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_0_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_0_2_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_0_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_1_0_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_1_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_1_1_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_1_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_1_2_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_1_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_2_0_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_2_0_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_2_1_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_2_1_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_I_2_2_t0b; // @[Top.scala 22:22]
  wire [7:0] n129_I_2_2_t1b; // @[Top.scala 22:22]
  wire [15:0] n129_O_0_0; // @[Top.scala 22:22]
  wire [15:0] n129_O_0_1; // @[Top.scala 22:22]
  wire [15:0] n129_O_0_2; // @[Top.scala 22:22]
  wire [15:0] n129_O_1_0; // @[Top.scala 22:22]
  wire [15:0] n129_O_1_1; // @[Top.scala 22:22]
  wire [15:0] n129_O_1_2; // @[Top.scala 22:22]
  wire [15:0] n129_O_2_0; // @[Top.scala 22:22]
  wire [15:0] n129_O_2_1; // @[Top.scala 22:22]
  wire [15:0] n129_O_2_2; // @[Top.scala 22:22]
  wire  n134_clock; // @[Top.scala 25:22]
  wire  n134_reset; // @[Top.scala 25:22]
  wire  n134_valid_up; // @[Top.scala 25:22]
  wire  n134_valid_down; // @[Top.scala 25:22]
  wire [15:0] n134_I_0_0; // @[Top.scala 25:22]
  wire [15:0] n134_I_0_1; // @[Top.scala 25:22]
  wire [15:0] n134_I_0_2; // @[Top.scala 25:22]
  wire [15:0] n134_I_1_0; // @[Top.scala 25:22]
  wire [15:0] n134_I_1_1; // @[Top.scala 25:22]
  wire [15:0] n134_I_1_2; // @[Top.scala 25:22]
  wire [15:0] n134_I_2_0; // @[Top.scala 25:22]
  wire [15:0] n134_I_2_1; // @[Top.scala 25:22]
  wire [15:0] n134_I_2_2; // @[Top.scala 25:22]
  wire [15:0] n134_O_0_0; // @[Top.scala 25:22]
  wire [15:0] n134_O_1_0; // @[Top.scala 25:22]
  wire [15:0] n134_O_2_0; // @[Top.scala 25:22]
  wire  n139_clock; // @[Top.scala 28:22]
  wire  n139_reset; // @[Top.scala 28:22]
  wire  n139_valid_up; // @[Top.scala 28:22]
  wire  n139_valid_down; // @[Top.scala 28:22]
  wire [15:0] n139_I_0_0; // @[Top.scala 28:22]
  wire [15:0] n139_I_1_0; // @[Top.scala 28:22]
  wire [15:0] n139_I_2_0; // @[Top.scala 28:22]
  wire [15:0] n139_O_0_0; // @[Top.scala 28:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n142_valid_up; // @[Top.scala 32:22]
  wire  n142_valid_down; // @[Top.scala 32:22]
  wire [15:0] n142_I0_0_0; // @[Top.scala 32:22]
  wire [15:0] n142_O_0_0_t0b; // @[Top.scala 32:22]
  wire [7:0] n142_O_0_0_t1b; // @[Top.scala 32:22]
  wire  n153_valid_up; // @[Top.scala 36:22]
  wire  n153_valid_down; // @[Top.scala 36:22]
  wire [15:0] n153_I_0_0_t0b; // @[Top.scala 36:22]
  wire [7:0] n153_I_0_0_t1b; // @[Top.scala 36:22]
  wire [15:0] n153_O_0_0; // @[Top.scala 36:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_9 n118 ( // @[Top.scala 18:22]
    .valid_up(n118_valid_up),
    .valid_down(n118_valid_down),
    .I0_0_0(n118_I0_0_0),
    .I0_0_1(n118_I0_0_1),
    .I0_0_2(n118_I0_0_2),
    .I0_1_0(n118_I0_1_0),
    .I0_1_1(n118_I0_1_1),
    .I0_1_2(n118_I0_1_2),
    .I0_2_0(n118_I0_2_0),
    .I0_2_1(n118_I0_2_1),
    .I0_2_2(n118_I0_2_2),
    .O_0_0_t0b(n118_O_0_0_t0b),
    .O_0_0_t1b(n118_O_0_0_t1b),
    .O_0_1_t0b(n118_O_0_1_t0b),
    .O_0_1_t1b(n118_O_0_1_t1b),
    .O_0_2_t0b(n118_O_0_2_t0b),
    .O_0_2_t1b(n118_O_0_2_t1b),
    .O_1_0_t0b(n118_O_1_0_t0b),
    .O_1_0_t1b(n118_O_1_0_t1b),
    .O_1_1_t0b(n118_O_1_1_t0b),
    .O_1_1_t1b(n118_O_1_1_t1b),
    .O_1_2_t0b(n118_O_1_2_t0b),
    .O_1_2_t1b(n118_O_1_2_t1b),
    .O_2_0_t0b(n118_O_2_0_t0b),
    .O_2_0_t1b(n118_O_2_0_t1b),
    .O_2_1_t0b(n118_O_2_1_t0b),
    .O_2_1_t1b(n118_O_2_1_t1b),
    .O_2_2_t0b(n118_O_2_2_t0b),
    .O_2_2_t1b(n118_O_2_2_t1b)
  );
  MapS_5 n129 ( // @[Top.scala 22:22]
    .valid_up(n129_valid_up),
    .valid_down(n129_valid_down),
    .I_0_0_t0b(n129_I_0_0_t0b),
    .I_0_0_t1b(n129_I_0_0_t1b),
    .I_0_1_t0b(n129_I_0_1_t0b),
    .I_0_1_t1b(n129_I_0_1_t1b),
    .I_0_2_t0b(n129_I_0_2_t0b),
    .I_0_2_t1b(n129_I_0_2_t1b),
    .I_1_0_t0b(n129_I_1_0_t0b),
    .I_1_0_t1b(n129_I_1_0_t1b),
    .I_1_1_t0b(n129_I_1_1_t0b),
    .I_1_1_t1b(n129_I_1_1_t1b),
    .I_1_2_t0b(n129_I_1_2_t0b),
    .I_1_2_t1b(n129_I_1_2_t1b),
    .I_2_0_t0b(n129_I_2_0_t0b),
    .I_2_0_t1b(n129_I_2_0_t1b),
    .I_2_1_t0b(n129_I_2_1_t0b),
    .I_2_1_t1b(n129_I_2_1_t1b),
    .I_2_2_t0b(n129_I_2_2_t0b),
    .I_2_2_t1b(n129_I_2_2_t1b),
    .O_0_0(n129_O_0_0),
    .O_0_1(n129_O_0_1),
    .O_0_2(n129_O_0_2),
    .O_1_0(n129_O_1_0),
    .O_1_1(n129_O_1_1),
    .O_1_2(n129_O_1_2),
    .O_2_0(n129_O_2_0),
    .O_2_1(n129_O_2_1),
    .O_2_2(n129_O_2_2)
  );
  MapS_6 n134 ( // @[Top.scala 25:22]
    .clock(n134_clock),
    .reset(n134_reset),
    .valid_up(n134_valid_up),
    .valid_down(n134_valid_down),
    .I_0_0(n134_I_0_0),
    .I_0_1(n134_I_0_1),
    .I_0_2(n134_I_0_2),
    .I_1_0(n134_I_1_0),
    .I_1_1(n134_I_1_1),
    .I_1_2(n134_I_1_2),
    .I_2_0(n134_I_2_0),
    .I_2_1(n134_I_2_1),
    .I_2_2(n134_I_2_2),
    .O_0_0(n134_O_0_0),
    .O_1_0(n134_O_1_0),
    .O_2_0(n134_O_2_0)
  );
  ReduceS_1 n139 ( // @[Top.scala 28:22]
    .clock(n139_clock),
    .reset(n139_reset),
    .valid_up(n139_valid_up),
    .valid_down(n139_valid_down),
    .I_0_0(n139_I_0_0),
    .I_1_0(n139_I_1_0),
    .I_2_0(n139_I_2_0),
    .O_0_0(n139_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n142 ( // @[Top.scala 32:22]
    .valid_up(n142_valid_up),
    .valid_down(n142_valid_down),
    .I0_0_0(n142_I0_0_0),
    .O_0_0_t0b(n142_O_0_0_t0b),
    .O_0_0_t1b(n142_O_0_0_t1b)
  );
  MapS_8 n153 ( // @[Top.scala 36:22]
    .valid_up(n153_valid_up),
    .valid_down(n153_valid_down),
    .I_0_0_t0b(n153_I_0_0_t0b),
    .I_0_0_t1b(n153_I_0_0_t1b),
    .O_0_0(n153_O_0_0)
  );
  assign valid_down = n153_valid_down; // @[Top.scala 40:16]
  assign O_0_0 = n153_O_0_0; // @[Top.scala 39:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n118_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 21:19]
  assign n118_I0_0_0 = I_0_0; // @[Top.scala 19:13]
  assign n118_I0_0_1 = I_0_1; // @[Top.scala 19:13]
  assign n118_I0_0_2 = I_0_2; // @[Top.scala 19:13]
  assign n118_I0_1_0 = I_1_0; // @[Top.scala 19:13]
  assign n118_I0_1_1 = I_1_1; // @[Top.scala 19:13]
  assign n118_I0_1_2 = I_1_2; // @[Top.scala 19:13]
  assign n118_I0_2_0 = I_2_0; // @[Top.scala 19:13]
  assign n118_I0_2_1 = I_2_1; // @[Top.scala 19:13]
  assign n118_I0_2_2 = I_2_2; // @[Top.scala 19:13]
  assign n129_valid_up = n118_valid_down; // @[Top.scala 24:19]
  assign n129_I_0_0_t0b = n118_O_0_0_t0b; // @[Top.scala 23:12]
  assign n129_I_0_0_t1b = n118_O_0_0_t1b; // @[Top.scala 23:12]
  assign n129_I_0_1_t0b = n118_O_0_1_t0b; // @[Top.scala 23:12]
  assign n129_I_0_1_t1b = n118_O_0_1_t1b; // @[Top.scala 23:12]
  assign n129_I_0_2_t0b = n118_O_0_2_t0b; // @[Top.scala 23:12]
  assign n129_I_0_2_t1b = n118_O_0_2_t1b; // @[Top.scala 23:12]
  assign n129_I_1_0_t0b = n118_O_1_0_t0b; // @[Top.scala 23:12]
  assign n129_I_1_0_t1b = n118_O_1_0_t1b; // @[Top.scala 23:12]
  assign n129_I_1_1_t0b = n118_O_1_1_t0b; // @[Top.scala 23:12]
  assign n129_I_1_1_t1b = n118_O_1_1_t1b; // @[Top.scala 23:12]
  assign n129_I_1_2_t0b = n118_O_1_2_t0b; // @[Top.scala 23:12]
  assign n129_I_1_2_t1b = n118_O_1_2_t1b; // @[Top.scala 23:12]
  assign n129_I_2_0_t0b = n118_O_2_0_t0b; // @[Top.scala 23:12]
  assign n129_I_2_0_t1b = n118_O_2_0_t1b; // @[Top.scala 23:12]
  assign n129_I_2_1_t0b = n118_O_2_1_t0b; // @[Top.scala 23:12]
  assign n129_I_2_1_t1b = n118_O_2_1_t1b; // @[Top.scala 23:12]
  assign n129_I_2_2_t0b = n118_O_2_2_t0b; // @[Top.scala 23:12]
  assign n129_I_2_2_t1b = n118_O_2_2_t1b; // @[Top.scala 23:12]
  assign n134_clock = clock;
  assign n134_reset = reset;
  assign n134_valid_up = n129_valid_down; // @[Top.scala 27:19]
  assign n134_I_0_0 = n129_O_0_0; // @[Top.scala 26:12]
  assign n134_I_0_1 = n129_O_0_1; // @[Top.scala 26:12]
  assign n134_I_0_2 = n129_O_0_2; // @[Top.scala 26:12]
  assign n134_I_1_0 = n129_O_1_0; // @[Top.scala 26:12]
  assign n134_I_1_1 = n129_O_1_1; // @[Top.scala 26:12]
  assign n134_I_1_2 = n129_O_1_2; // @[Top.scala 26:12]
  assign n134_I_2_0 = n129_O_2_0; // @[Top.scala 26:12]
  assign n134_I_2_1 = n129_O_2_1; // @[Top.scala 26:12]
  assign n134_I_2_2 = n129_O_2_2; // @[Top.scala 26:12]
  assign n139_clock = clock;
  assign n139_reset = reset;
  assign n139_valid_up = n134_valid_down; // @[Top.scala 30:19]
  assign n139_I_0_0 = n134_O_0_0; // @[Top.scala 29:12]
  assign n139_I_1_0 = n134_O_1_0; // @[Top.scala 29:12]
  assign n139_I_2_0 = n134_O_2_0; // @[Top.scala 29:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n142_valid_up = n139_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 35:19]
  assign n142_I0_0_0 = n139_O_0_0; // @[Top.scala 33:13]
  assign n153_valid_up = n142_valid_down; // @[Top.scala 38:19]
  assign n153_I_0_0_t0b = n142_O_0_0_t0b; // @[Top.scala 37:12]
  assign n153_I_0_0_t1b = n142_O_0_0_t1b; // @[Top.scala 37:12]
endmodule
module MapS_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  input  [15:0] I_8_0_0,
  input  [15:0] I_8_0_1,
  input  [15:0] I_8_0_2,
  input  [15:0] I_8_1_0,
  input  [15:0] I_8_1_1,
  input  [15:0] I_8_1_2,
  input  [15:0] I_8_2_0,
  input  [15:0] I_8_2_1,
  input  [15:0] I_8_2_2,
  input  [15:0] I_9_0_0,
  input  [15:0] I_9_0_1,
  input  [15:0] I_9_0_2,
  input  [15:0] I_9_1_0,
  input  [15:0] I_9_1_1,
  input  [15:0] I_9_1_2,
  input  [15:0] I_9_2_0,
  input  [15:0] I_9_2_1,
  input  [15:0] I_9_2_2,
  input  [15:0] I_10_0_0,
  input  [15:0] I_10_0_1,
  input  [15:0] I_10_0_2,
  input  [15:0] I_10_1_0,
  input  [15:0] I_10_1_1,
  input  [15:0] I_10_1_2,
  input  [15:0] I_10_2_0,
  input  [15:0] I_10_2_1,
  input  [15:0] I_10_2_2,
  input  [15:0] I_11_0_0,
  input  [15:0] I_11_0_1,
  input  [15:0] I_11_0_2,
  input  [15:0] I_11_1_0,
  input  [15:0] I_11_1_1,
  input  [15:0] I_11_1_2,
  input  [15:0] I_11_2_0,
  input  [15:0] I_11_2_1,
  input  [15:0] I_11_2_2,
  input  [15:0] I_12_0_0,
  input  [15:0] I_12_0_1,
  input  [15:0] I_12_0_2,
  input  [15:0] I_12_1_0,
  input  [15:0] I_12_1_1,
  input  [15:0] I_12_1_2,
  input  [15:0] I_12_2_0,
  input  [15:0] I_12_2_1,
  input  [15:0] I_12_2_2,
  input  [15:0] I_13_0_0,
  input  [15:0] I_13_0_1,
  input  [15:0] I_13_0_2,
  input  [15:0] I_13_1_0,
  input  [15:0] I_13_1_1,
  input  [15:0] I_13_1_2,
  input  [15:0] I_13_2_0,
  input  [15:0] I_13_2_1,
  input  [15:0] I_13_2_2,
  input  [15:0] I_14_0_0,
  input  [15:0] I_14_0_1,
  input  [15:0] I_14_0_2,
  input  [15:0] I_14_1_0,
  input  [15:0] I_14_1_1,
  input  [15:0] I_14_1_2,
  input  [15:0] I_14_2_0,
  input  [15:0] I_14_2_1,
  input  [15:0] I_14_2_2,
  input  [15:0] I_15_0_0,
  input  [15:0] I_15_0_1,
  input  [15:0] I_15_0_2,
  input  [15:0] I_15_1_0,
  input  [15:0] I_15_1_1,
  input  [15:0] I_15_1_2,
  input  [15:0] I_15_2_0,
  input  [15:0] I_15_2_1,
  input  [15:0] I_15_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0,
  output [15:0] O_4_0_0,
  output [15:0] O_5_0_0,
  output [15:0] O_6_0_0,
  output [15:0] O_7_0_0,
  output [15:0] O_8_0_0,
  output [15:0] O_9_0_0,
  output [15:0] O_10_0_0,
  output [15:0] O_11_0_0,
  output [15:0] O_12_0_0,
  output [15:0] O_13_0_0,
  output [15:0] O_14_0_0,
  output [15:0] O_15_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [15:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [15:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_7_clock; // @[MapS.scala 10:86]
  wire  other_ops_7_reset; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_8_clock; // @[MapS.scala 10:86]
  wire  other_ops_8_reset; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_9_clock; // @[MapS.scala 10:86]
  wire  other_ops_9_reset; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_10_clock; // @[MapS.scala 10:86]
  wire  other_ops_10_reset; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_11_clock; // @[MapS.scala 10:86]
  wire  other_ops_11_reset; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_12_clock; // @[MapS.scala 10:86]
  wire  other_ops_12_reset; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_13_clock; // @[MapS.scala 10:86]
  wire  other_ops_13_reset; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_14_clock; // @[MapS.scala 10:86]
  wire  other_ops_14_reset; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_1_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_1_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_1_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_2_0; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_2_1; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_I_2_2; // @[MapS.scala 10:86]
  wire [15:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  Module_0 other_ops_7 ( // @[MapS.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .I_1_0(other_ops_7_I_1_0),
    .I_1_1(other_ops_7_I_1_1),
    .I_1_2(other_ops_7_I_1_2),
    .I_2_0(other_ops_7_I_2_0),
    .I_2_1(other_ops_7_I_2_1),
    .I_2_2(other_ops_7_I_2_2),
    .O_0_0(other_ops_7_O_0_0)
  );
  Module_0 other_ops_8 ( // @[MapS.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .I_1_0(other_ops_8_I_1_0),
    .I_1_1(other_ops_8_I_1_1),
    .I_1_2(other_ops_8_I_1_2),
    .I_2_0(other_ops_8_I_2_0),
    .I_2_1(other_ops_8_I_2_1),
    .I_2_2(other_ops_8_I_2_2),
    .O_0_0(other_ops_8_O_0_0)
  );
  Module_0 other_ops_9 ( // @[MapS.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .I_1_0(other_ops_9_I_1_0),
    .I_1_1(other_ops_9_I_1_1),
    .I_1_2(other_ops_9_I_1_2),
    .I_2_0(other_ops_9_I_2_0),
    .I_2_1(other_ops_9_I_2_1),
    .I_2_2(other_ops_9_I_2_2),
    .O_0_0(other_ops_9_O_0_0)
  );
  Module_0 other_ops_10 ( // @[MapS.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .I_1_0(other_ops_10_I_1_0),
    .I_1_1(other_ops_10_I_1_1),
    .I_1_2(other_ops_10_I_1_2),
    .I_2_0(other_ops_10_I_2_0),
    .I_2_1(other_ops_10_I_2_1),
    .I_2_2(other_ops_10_I_2_2),
    .O_0_0(other_ops_10_O_0_0)
  );
  Module_0 other_ops_11 ( // @[MapS.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .I_1_0(other_ops_11_I_1_0),
    .I_1_1(other_ops_11_I_1_1),
    .I_1_2(other_ops_11_I_1_2),
    .I_2_0(other_ops_11_I_2_0),
    .I_2_1(other_ops_11_I_2_1),
    .I_2_2(other_ops_11_I_2_2),
    .O_0_0(other_ops_11_O_0_0)
  );
  Module_0 other_ops_12 ( // @[MapS.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .I_1_0(other_ops_12_I_1_0),
    .I_1_1(other_ops_12_I_1_1),
    .I_1_2(other_ops_12_I_1_2),
    .I_2_0(other_ops_12_I_2_0),
    .I_2_1(other_ops_12_I_2_1),
    .I_2_2(other_ops_12_I_2_2),
    .O_0_0(other_ops_12_O_0_0)
  );
  Module_0 other_ops_13 ( // @[MapS.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .I_1_0(other_ops_13_I_1_0),
    .I_1_1(other_ops_13_I_1_1),
    .I_1_2(other_ops_13_I_1_2),
    .I_2_0(other_ops_13_I_2_0),
    .I_2_1(other_ops_13_I_2_1),
    .I_2_2(other_ops_13_I_2_2),
    .O_0_0(other_ops_13_O_0_0)
  );
  Module_0 other_ops_14 ( // @[MapS.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .I_1_0(other_ops_14_I_1_0),
    .I_1_1(other_ops_14_I_1_1),
    .I_1_2(other_ops_14_I_1_2),
    .I_2_0(other_ops_14_I_2_0),
    .I_2_1(other_ops_14_I_2_1),
    .I_2_2(other_ops_14_I_2_2),
    .O_0_0(other_ops_14_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_7_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_0 = I_8_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_1 = I_8_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_2 = I_8_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_0 = I_8_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_1 = I_8_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_2 = I_8_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_8_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_0 = I_9_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_1 = I_9_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_2 = I_9_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_0 = I_9_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_1 = I_9_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_2 = I_9_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_9_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_0 = I_10_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_1 = I_10_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_2 = I_10_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_0 = I_10_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_1 = I_10_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_2 = I_10_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_10_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_0 = I_11_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_1 = I_11_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_2 = I_11_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_0 = I_11_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_1 = I_11_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_2 = I_11_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_11_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_0 = I_12_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_1 = I_12_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_2 = I_12_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_0 = I_12_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_1 = I_12_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_2 = I_12_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_12_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_0 = I_13_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_1 = I_13_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_2 = I_13_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_0 = I_13_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_1 = I_13_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_2 = I_13_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_13_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_0 = I_14_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_1 = I_14_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_2 = I_14_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_0 = I_14_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_1 = I_14_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_2 = I_14_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_14_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_0 = I_15_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_1 = I_15_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_2 = I_15_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_0 = I_15_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_1 = I_15_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_2 = I_15_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_8(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_0_0_1,
  input  [15:0] I_0_0_2,
  input  [15:0] I_0_1_0,
  input  [15:0] I_0_1_1,
  input  [15:0] I_0_1_2,
  input  [15:0] I_0_2_0,
  input  [15:0] I_0_2_1,
  input  [15:0] I_0_2_2,
  input  [15:0] I_1_0_0,
  input  [15:0] I_1_0_1,
  input  [15:0] I_1_0_2,
  input  [15:0] I_1_1_0,
  input  [15:0] I_1_1_1,
  input  [15:0] I_1_1_2,
  input  [15:0] I_1_2_0,
  input  [15:0] I_1_2_1,
  input  [15:0] I_1_2_2,
  input  [15:0] I_2_0_0,
  input  [15:0] I_2_0_1,
  input  [15:0] I_2_0_2,
  input  [15:0] I_2_1_0,
  input  [15:0] I_2_1_1,
  input  [15:0] I_2_1_2,
  input  [15:0] I_2_2_0,
  input  [15:0] I_2_2_1,
  input  [15:0] I_2_2_2,
  input  [15:0] I_3_0_0,
  input  [15:0] I_3_0_1,
  input  [15:0] I_3_0_2,
  input  [15:0] I_3_1_0,
  input  [15:0] I_3_1_1,
  input  [15:0] I_3_1_2,
  input  [15:0] I_3_2_0,
  input  [15:0] I_3_2_1,
  input  [15:0] I_3_2_2,
  input  [15:0] I_4_0_0,
  input  [15:0] I_4_0_1,
  input  [15:0] I_4_0_2,
  input  [15:0] I_4_1_0,
  input  [15:0] I_4_1_1,
  input  [15:0] I_4_1_2,
  input  [15:0] I_4_2_0,
  input  [15:0] I_4_2_1,
  input  [15:0] I_4_2_2,
  input  [15:0] I_5_0_0,
  input  [15:0] I_5_0_1,
  input  [15:0] I_5_0_2,
  input  [15:0] I_5_1_0,
  input  [15:0] I_5_1_1,
  input  [15:0] I_5_1_2,
  input  [15:0] I_5_2_0,
  input  [15:0] I_5_2_1,
  input  [15:0] I_5_2_2,
  input  [15:0] I_6_0_0,
  input  [15:0] I_6_0_1,
  input  [15:0] I_6_0_2,
  input  [15:0] I_6_1_0,
  input  [15:0] I_6_1_1,
  input  [15:0] I_6_1_2,
  input  [15:0] I_6_2_0,
  input  [15:0] I_6_2_1,
  input  [15:0] I_6_2_2,
  input  [15:0] I_7_0_0,
  input  [15:0] I_7_0_1,
  input  [15:0] I_7_0_2,
  input  [15:0] I_7_1_0,
  input  [15:0] I_7_1_1,
  input  [15:0] I_7_1_2,
  input  [15:0] I_7_2_0,
  input  [15:0] I_7_2_1,
  input  [15:0] I_7_2_2,
  input  [15:0] I_8_0_0,
  input  [15:0] I_8_0_1,
  input  [15:0] I_8_0_2,
  input  [15:0] I_8_1_0,
  input  [15:0] I_8_1_1,
  input  [15:0] I_8_1_2,
  input  [15:0] I_8_2_0,
  input  [15:0] I_8_2_1,
  input  [15:0] I_8_2_2,
  input  [15:0] I_9_0_0,
  input  [15:0] I_9_0_1,
  input  [15:0] I_9_0_2,
  input  [15:0] I_9_1_0,
  input  [15:0] I_9_1_1,
  input  [15:0] I_9_1_2,
  input  [15:0] I_9_2_0,
  input  [15:0] I_9_2_1,
  input  [15:0] I_9_2_2,
  input  [15:0] I_10_0_0,
  input  [15:0] I_10_0_1,
  input  [15:0] I_10_0_2,
  input  [15:0] I_10_1_0,
  input  [15:0] I_10_1_1,
  input  [15:0] I_10_1_2,
  input  [15:0] I_10_2_0,
  input  [15:0] I_10_2_1,
  input  [15:0] I_10_2_2,
  input  [15:0] I_11_0_0,
  input  [15:0] I_11_0_1,
  input  [15:0] I_11_0_2,
  input  [15:0] I_11_1_0,
  input  [15:0] I_11_1_1,
  input  [15:0] I_11_1_2,
  input  [15:0] I_11_2_0,
  input  [15:0] I_11_2_1,
  input  [15:0] I_11_2_2,
  input  [15:0] I_12_0_0,
  input  [15:0] I_12_0_1,
  input  [15:0] I_12_0_2,
  input  [15:0] I_12_1_0,
  input  [15:0] I_12_1_1,
  input  [15:0] I_12_1_2,
  input  [15:0] I_12_2_0,
  input  [15:0] I_12_2_1,
  input  [15:0] I_12_2_2,
  input  [15:0] I_13_0_0,
  input  [15:0] I_13_0_1,
  input  [15:0] I_13_0_2,
  input  [15:0] I_13_1_0,
  input  [15:0] I_13_1_1,
  input  [15:0] I_13_1_2,
  input  [15:0] I_13_2_0,
  input  [15:0] I_13_2_1,
  input  [15:0] I_13_2_2,
  input  [15:0] I_14_0_0,
  input  [15:0] I_14_0_1,
  input  [15:0] I_14_0_2,
  input  [15:0] I_14_1_0,
  input  [15:0] I_14_1_1,
  input  [15:0] I_14_1_2,
  input  [15:0] I_14_2_0,
  input  [15:0] I_14_2_1,
  input  [15:0] I_14_2_2,
  input  [15:0] I_15_0_0,
  input  [15:0] I_15_0_1,
  input  [15:0] I_15_0_2,
  input  [15:0] I_15_1_0,
  input  [15:0] I_15_1_1,
  input  [15:0] I_15_1_2,
  input  [15:0] I_15_2_0,
  input  [15:0] I_15_2_1,
  input  [15:0] I_15_2_2,
  output [15:0] O_0_0_0,
  output [15:0] O_1_0_0,
  output [15:0] O_2_0_0,
  output [15:0] O_3_0_0,
  output [15:0] O_4_0_0,
  output [15:0] O_5_0_0,
  output [15:0] O_6_0_0,
  output [15:0] O_7_0_0,
  output [15:0] O_8_0_0,
  output [15:0] O_9_0_0,
  output [15:0] O_10_0_0,
  output [15:0] O_11_0_0,
  output [15:0] O_12_0_0,
  output [15:0] O_13_0_0,
  output [15:0] O_14_0_0,
  output [15:0] O_15_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_8_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_9_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_10_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_11_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_12_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_13_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_14_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_1_2; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_2_0; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_2_1; // @[MapT.scala 8:20]
  wire [15:0] op_I_15_2_2; // @[MapT.scala 8:20]
  wire [15:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [15:0] op_O_15_0_0; // @[MapT.scala 8:20]
  MapS_9 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_8_1_2(op_I_8_1_2),
    .I_8_2_0(op_I_8_2_0),
    .I_8_2_1(op_I_8_2_1),
    .I_8_2_2(op_I_8_2_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_9_1_2(op_I_9_1_2),
    .I_9_2_0(op_I_9_2_0),
    .I_9_2_1(op_I_9_2_1),
    .I_9_2_2(op_I_9_2_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_10_1_2(op_I_10_1_2),
    .I_10_2_0(op_I_10_2_0),
    .I_10_2_1(op_I_10_2_1),
    .I_10_2_2(op_I_10_2_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_11_1_2(op_I_11_1_2),
    .I_11_2_0(op_I_11_2_0),
    .I_11_2_1(op_I_11_2_1),
    .I_11_2_2(op_I_11_2_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_12_1_2(op_I_12_1_2),
    .I_12_2_0(op_I_12_2_0),
    .I_12_2_1(op_I_12_2_1),
    .I_12_2_2(op_I_12_2_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_13_1_2(op_I_13_1_2),
    .I_13_2_0(op_I_13_2_0),
    .I_13_2_1(op_I_13_2_1),
    .I_13_2_2(op_I_13_2_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_14_1_2(op_I_14_1_2),
    .I_14_2_0(op_I_14_2_0),
    .I_14_2_1(op_I_14_2_1),
    .I_14_2_2(op_I_14_2_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .I_15_1_2(op_I_15_1_2),
    .I_15_2_0(op_I_15_2_0),
    .I_15_2_1(op_I_15_2_1),
    .I_15_2_2(op_I_15_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0),
    .O_8_0_0(op_O_8_0_0),
    .O_9_0_0(op_O_9_0_0),
    .O_10_0_0(op_O_10_0_0),
    .O_11_0_0(op_O_11_0_0),
    .O_12_0_0(op_O_12_0_0),
    .O_13_0_0(op_O_13_0_0),
    .O_14_0_0(op_O_14_0_0),
    .O_15_0_0(op_O_15_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_8_1_2 = I_8_1_2; // @[MapT.scala 14:10]
  assign op_I_8_2_0 = I_8_2_0; // @[MapT.scala 14:10]
  assign op_I_8_2_1 = I_8_2_1; // @[MapT.scala 14:10]
  assign op_I_8_2_2 = I_8_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_9_1_2 = I_9_1_2; // @[MapT.scala 14:10]
  assign op_I_9_2_0 = I_9_2_0; // @[MapT.scala 14:10]
  assign op_I_9_2_1 = I_9_2_1; // @[MapT.scala 14:10]
  assign op_I_9_2_2 = I_9_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_10_1_2 = I_10_1_2; // @[MapT.scala 14:10]
  assign op_I_10_2_0 = I_10_2_0; // @[MapT.scala 14:10]
  assign op_I_10_2_1 = I_10_2_1; // @[MapT.scala 14:10]
  assign op_I_10_2_2 = I_10_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_11_1_2 = I_11_1_2; // @[MapT.scala 14:10]
  assign op_I_11_2_0 = I_11_2_0; // @[MapT.scala 14:10]
  assign op_I_11_2_1 = I_11_2_1; // @[MapT.scala 14:10]
  assign op_I_11_2_2 = I_11_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_12_1_2 = I_12_1_2; // @[MapT.scala 14:10]
  assign op_I_12_2_0 = I_12_2_0; // @[MapT.scala 14:10]
  assign op_I_12_2_1 = I_12_2_1; // @[MapT.scala 14:10]
  assign op_I_12_2_2 = I_12_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_13_1_2 = I_13_1_2; // @[MapT.scala 14:10]
  assign op_I_13_2_0 = I_13_2_0; // @[MapT.scala 14:10]
  assign op_I_13_2_1 = I_13_2_1; // @[MapT.scala 14:10]
  assign op_I_13_2_2 = I_13_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_14_1_2 = I_14_1_2; // @[MapT.scala 14:10]
  assign op_I_14_2_0 = I_14_2_0; // @[MapT.scala 14:10]
  assign op_I_14_2_1 = I_14_2_1; // @[MapT.scala 14:10]
  assign op_I_14_2_2 = I_14_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
  assign op_I_15_1_2 = I_15_1_2; // @[MapT.scala 14:10]
  assign op_I_15_2_0 = I_15_2_0; // @[MapT.scala 14:10]
  assign op_I_15_2_1 = I_15_2_1; // @[MapT.scala 14:10]
  assign op_I_15_2_2 = I_15_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0_0,
  input  [15:0] I_1_0_0,
  input  [15:0] I_2_0_0,
  input  [15:0] I_3_0_0,
  input  [15:0] I_4_0_0,
  input  [15:0] I_5_0_0,
  input  [15:0] I_6_0_0,
  input  [15:0] I_7_0_0,
  input  [15:0] I_8_0_0,
  input  [15:0] I_9_0_0,
  input  [15:0] I_10_0_0,
  input  [15:0] I_11_0_0,
  input  [15:0] I_12_0_0,
  input  [15:0] I_13_0_0,
  input  [15:0] I_14_0_0,
  input  [15:0] I_15_0_0,
  output [15:0] O_0_0,
  output [15:0] O_1_0,
  output [15:0] O_2_0,
  output [15:0] O_3_0,
  output [15:0] O_4_0,
  output [15:0] O_5_0,
  output [15:0] O_6_0,
  output [15:0] O_7_0,
  output [15:0] O_8_0,
  output [15:0] O_9_0,
  output [15:0] O_10_0,
  output [15:0] O_11_0,
  output [15:0] O_12_0,
  output [15:0] O_13_0,
  output [15:0] O_14_0,
  output [15:0] O_15_0
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0 = I_1_0_0; // @[Passthrough.scala 17:68]
  assign O_2_0 = I_2_0_0; // @[Passthrough.scala 17:68]
  assign O_3_0 = I_3_0_0; // @[Passthrough.scala 17:68]
  assign O_4_0 = I_4_0_0; // @[Passthrough.scala 17:68]
  assign O_5_0 = I_5_0_0; // @[Passthrough.scala 17:68]
  assign O_6_0 = I_6_0_0; // @[Passthrough.scala 17:68]
  assign O_7_0 = I_7_0_0; // @[Passthrough.scala 17:68]
  assign O_8_0 = I_8_0_0; // @[Passthrough.scala 17:68]
  assign O_9_0 = I_9_0_0; // @[Passthrough.scala 17:68]
  assign O_10_0 = I_10_0_0; // @[Passthrough.scala 17:68]
  assign O_11_0 = I_11_0_0; // @[Passthrough.scala 17:68]
  assign O_12_0 = I_12_0_0; // @[Passthrough.scala 17:68]
  assign O_13_0 = I_13_0_0; // @[Passthrough.scala 17:68]
  assign O_14_0 = I_14_0_0; // @[Passthrough.scala 17:68]
  assign O_15_0 = I_15_0_0; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_1(
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0_0,
  input  [15:0] I_1_0,
  input  [15:0] I_2_0,
  input  [15:0] I_3_0,
  input  [15:0] I_4_0,
  input  [15:0] I_5_0,
  input  [15:0] I_6_0,
  input  [15:0] I_7_0,
  input  [15:0] I_8_0,
  input  [15:0] I_9_0,
  input  [15:0] I_10_0,
  input  [15:0] I_11_0,
  input  [15:0] I_12_0,
  input  [15:0] I_13_0,
  input  [15:0] I_14_0,
  input  [15:0] I_15_0,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7,
  output [15:0] O_8,
  output [15:0] O_9,
  output [15:0] O_10,
  output [15:0] O_11,
  output [15:0] O_12,
  output [15:0] O_13,
  output [15:0] O_14,
  output [15:0] O_15
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_1_0; // @[Passthrough.scala 17:68]
  assign O_2 = I_2_0; // @[Passthrough.scala 17:68]
  assign O_3 = I_3_0; // @[Passthrough.scala 17:68]
  assign O_4 = I_4_0; // @[Passthrough.scala 17:68]
  assign O_5 = I_5_0; // @[Passthrough.scala 17:68]
  assign O_6 = I_6_0; // @[Passthrough.scala 17:68]
  assign O_7 = I_7_0; // @[Passthrough.scala 17:68]
  assign O_8 = I_8_0; // @[Passthrough.scala 17:68]
  assign O_9 = I_9_0; // @[Passthrough.scala 17:68]
  assign O_10 = I_10_0; // @[Passthrough.scala 17:68]
  assign O_11 = I_11_0; // @[Passthrough.scala 17:68]
  assign O_12 = I_12_0; // @[Passthrough.scala 17:68]
  assign O_13 = I_13_0; // @[Passthrough.scala 17:68]
  assign O_14 = I_14_0; // @[Passthrough.scala 17:68]
  assign O_15 = I_15_0; // @[Passthrough.scala 17:68]
endmodule
module Top(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [15:0] I_0,
  input  [15:0] I_1,
  input  [15:0] I_2,
  input  [15:0] I_3,
  input  [15:0] I_4,
  input  [15:0] I_5,
  input  [15:0] I_6,
  input  [15:0] I_7,
  input  [15:0] I_8,
  input  [15:0] I_9,
  input  [15:0] I_10,
  input  [15:0] I_11,
  input  [15:0] I_12,
  input  [15:0] I_13,
  input  [15:0] I_14,
  input  [15:0] I_15,
  output [15:0] O_0,
  output [15:0] O_1,
  output [15:0] O_2,
  output [15:0] O_3,
  output [15:0] O_4,
  output [15:0] O_5,
  output [15:0] O_6,
  output [15:0] O_7,
  output [15:0] O_8,
  output [15:0] O_9,
  output [15:0] O_10,
  output [15:0] O_11,
  output [15:0] O_12,
  output [15:0] O_13,
  output [15:0] O_14,
  output [15:0] O_15
);
  wire  n1_clock; // @[Top.scala 46:20]
  wire  n1_reset; // @[Top.scala 46:20]
  wire  n1_valid_up; // @[Top.scala 46:20]
  wire  n1_valid_down; // @[Top.scala 46:20]
  wire [15:0] n1_I_0; // @[Top.scala 46:20]
  wire [15:0] n1_I_1; // @[Top.scala 46:20]
  wire [15:0] n1_I_2; // @[Top.scala 46:20]
  wire [15:0] n1_I_3; // @[Top.scala 46:20]
  wire [15:0] n1_I_4; // @[Top.scala 46:20]
  wire [15:0] n1_I_5; // @[Top.scala 46:20]
  wire [15:0] n1_I_6; // @[Top.scala 46:20]
  wire [15:0] n1_I_7; // @[Top.scala 46:20]
  wire [15:0] n1_I_8; // @[Top.scala 46:20]
  wire [15:0] n1_I_9; // @[Top.scala 46:20]
  wire [15:0] n1_I_10; // @[Top.scala 46:20]
  wire [15:0] n1_I_11; // @[Top.scala 46:20]
  wire [15:0] n1_I_12; // @[Top.scala 46:20]
  wire [15:0] n1_I_13; // @[Top.scala 46:20]
  wire [15:0] n1_I_14; // @[Top.scala 46:20]
  wire [15:0] n1_I_15; // @[Top.scala 46:20]
  wire [15:0] n1_O_0; // @[Top.scala 46:20]
  wire [15:0] n1_O_1; // @[Top.scala 46:20]
  wire [15:0] n1_O_2; // @[Top.scala 46:20]
  wire [15:0] n1_O_3; // @[Top.scala 46:20]
  wire [15:0] n1_O_4; // @[Top.scala 46:20]
  wire [15:0] n1_O_5; // @[Top.scala 46:20]
  wire [15:0] n1_O_6; // @[Top.scala 46:20]
  wire [15:0] n1_O_7; // @[Top.scala 46:20]
  wire [15:0] n1_O_8; // @[Top.scala 46:20]
  wire [15:0] n1_O_9; // @[Top.scala 46:20]
  wire [15:0] n1_O_10; // @[Top.scala 46:20]
  wire [15:0] n1_O_11; // @[Top.scala 46:20]
  wire [15:0] n1_O_12; // @[Top.scala 46:20]
  wire [15:0] n1_O_13; // @[Top.scala 46:20]
  wire [15:0] n1_O_14; // @[Top.scala 46:20]
  wire [15:0] n1_O_15; // @[Top.scala 46:20]
  wire  n2_clock; // @[Top.scala 49:20]
  wire  n2_reset; // @[Top.scala 49:20]
  wire  n2_valid_up; // @[Top.scala 49:20]
  wire  n2_valid_down; // @[Top.scala 49:20]
  wire [15:0] n2_I_0; // @[Top.scala 49:20]
  wire [15:0] n2_I_1; // @[Top.scala 49:20]
  wire [15:0] n2_I_2; // @[Top.scala 49:20]
  wire [15:0] n2_I_3; // @[Top.scala 49:20]
  wire [15:0] n2_I_4; // @[Top.scala 49:20]
  wire [15:0] n2_I_5; // @[Top.scala 49:20]
  wire [15:0] n2_I_6; // @[Top.scala 49:20]
  wire [15:0] n2_I_7; // @[Top.scala 49:20]
  wire [15:0] n2_I_8; // @[Top.scala 49:20]
  wire [15:0] n2_I_9; // @[Top.scala 49:20]
  wire [15:0] n2_I_10; // @[Top.scala 49:20]
  wire [15:0] n2_I_11; // @[Top.scala 49:20]
  wire [15:0] n2_I_12; // @[Top.scala 49:20]
  wire [15:0] n2_I_13; // @[Top.scala 49:20]
  wire [15:0] n2_I_14; // @[Top.scala 49:20]
  wire [15:0] n2_I_15; // @[Top.scala 49:20]
  wire [15:0] n2_O_0; // @[Top.scala 49:20]
  wire [15:0] n2_O_1; // @[Top.scala 49:20]
  wire [15:0] n2_O_2; // @[Top.scala 49:20]
  wire [15:0] n2_O_3; // @[Top.scala 49:20]
  wire [15:0] n2_O_4; // @[Top.scala 49:20]
  wire [15:0] n2_O_5; // @[Top.scala 49:20]
  wire [15:0] n2_O_6; // @[Top.scala 49:20]
  wire [15:0] n2_O_7; // @[Top.scala 49:20]
  wire [15:0] n2_O_8; // @[Top.scala 49:20]
  wire [15:0] n2_O_9; // @[Top.scala 49:20]
  wire [15:0] n2_O_10; // @[Top.scala 49:20]
  wire [15:0] n2_O_11; // @[Top.scala 49:20]
  wire [15:0] n2_O_12; // @[Top.scala 49:20]
  wire [15:0] n2_O_13; // @[Top.scala 49:20]
  wire [15:0] n2_O_14; // @[Top.scala 49:20]
  wire [15:0] n2_O_15; // @[Top.scala 49:20]
  wire  n3_clock; // @[Top.scala 52:20]
  wire  n3_reset; // @[Top.scala 52:20]
  wire  n3_valid_up; // @[Top.scala 52:20]
  wire  n3_valid_down; // @[Top.scala 52:20]
  wire [15:0] n3_I_0; // @[Top.scala 52:20]
  wire [15:0] n3_I_1; // @[Top.scala 52:20]
  wire [15:0] n3_I_2; // @[Top.scala 52:20]
  wire [15:0] n3_I_3; // @[Top.scala 52:20]
  wire [15:0] n3_I_4; // @[Top.scala 52:20]
  wire [15:0] n3_I_5; // @[Top.scala 52:20]
  wire [15:0] n3_I_6; // @[Top.scala 52:20]
  wire [15:0] n3_I_7; // @[Top.scala 52:20]
  wire [15:0] n3_I_8; // @[Top.scala 52:20]
  wire [15:0] n3_I_9; // @[Top.scala 52:20]
  wire [15:0] n3_I_10; // @[Top.scala 52:20]
  wire [15:0] n3_I_11; // @[Top.scala 52:20]
  wire [15:0] n3_I_12; // @[Top.scala 52:20]
  wire [15:0] n3_I_13; // @[Top.scala 52:20]
  wire [15:0] n3_I_14; // @[Top.scala 52:20]
  wire [15:0] n3_I_15; // @[Top.scala 52:20]
  wire [15:0] n3_O_0; // @[Top.scala 52:20]
  wire [15:0] n3_O_1; // @[Top.scala 52:20]
  wire [15:0] n3_O_2; // @[Top.scala 52:20]
  wire [15:0] n3_O_3; // @[Top.scala 52:20]
  wire [15:0] n3_O_4; // @[Top.scala 52:20]
  wire [15:0] n3_O_5; // @[Top.scala 52:20]
  wire [15:0] n3_O_6; // @[Top.scala 52:20]
  wire [15:0] n3_O_7; // @[Top.scala 52:20]
  wire [15:0] n3_O_8; // @[Top.scala 52:20]
  wire [15:0] n3_O_9; // @[Top.scala 52:20]
  wire [15:0] n3_O_10; // @[Top.scala 52:20]
  wire [15:0] n3_O_11; // @[Top.scala 52:20]
  wire [15:0] n3_O_12; // @[Top.scala 52:20]
  wire [15:0] n3_O_13; // @[Top.scala 52:20]
  wire [15:0] n3_O_14; // @[Top.scala 52:20]
  wire [15:0] n3_O_15; // @[Top.scala 52:20]
  wire  n4_clock; // @[Top.scala 55:20]
  wire  n4_reset; // @[Top.scala 55:20]
  wire  n4_valid_up; // @[Top.scala 55:20]
  wire  n4_valid_down; // @[Top.scala 55:20]
  wire [15:0] n4_I_0; // @[Top.scala 55:20]
  wire [15:0] n4_I_1; // @[Top.scala 55:20]
  wire [15:0] n4_I_2; // @[Top.scala 55:20]
  wire [15:0] n4_I_3; // @[Top.scala 55:20]
  wire [15:0] n4_I_4; // @[Top.scala 55:20]
  wire [15:0] n4_I_5; // @[Top.scala 55:20]
  wire [15:0] n4_I_6; // @[Top.scala 55:20]
  wire [15:0] n4_I_7; // @[Top.scala 55:20]
  wire [15:0] n4_I_8; // @[Top.scala 55:20]
  wire [15:0] n4_I_9; // @[Top.scala 55:20]
  wire [15:0] n4_I_10; // @[Top.scala 55:20]
  wire [15:0] n4_I_11; // @[Top.scala 55:20]
  wire [15:0] n4_I_12; // @[Top.scala 55:20]
  wire [15:0] n4_I_13; // @[Top.scala 55:20]
  wire [15:0] n4_I_14; // @[Top.scala 55:20]
  wire [15:0] n4_I_15; // @[Top.scala 55:20]
  wire [15:0] n4_O_0; // @[Top.scala 55:20]
  wire [15:0] n4_O_1; // @[Top.scala 55:20]
  wire [15:0] n4_O_2; // @[Top.scala 55:20]
  wire [15:0] n4_O_3; // @[Top.scala 55:20]
  wire [15:0] n4_O_4; // @[Top.scala 55:20]
  wire [15:0] n4_O_5; // @[Top.scala 55:20]
  wire [15:0] n4_O_6; // @[Top.scala 55:20]
  wire [15:0] n4_O_7; // @[Top.scala 55:20]
  wire [15:0] n4_O_8; // @[Top.scala 55:20]
  wire [15:0] n4_O_9; // @[Top.scala 55:20]
  wire [15:0] n4_O_10; // @[Top.scala 55:20]
  wire [15:0] n4_O_11; // @[Top.scala 55:20]
  wire [15:0] n4_O_12; // @[Top.scala 55:20]
  wire [15:0] n4_O_13; // @[Top.scala 55:20]
  wire [15:0] n4_O_14; // @[Top.scala 55:20]
  wire [15:0] n4_O_15; // @[Top.scala 55:20]
  wire  n5_clock; // @[Top.scala 58:20]
  wire  n5_reset; // @[Top.scala 58:20]
  wire  n5_valid_up; // @[Top.scala 58:20]
  wire  n5_valid_down; // @[Top.scala 58:20]
  wire [15:0] n5_I_0; // @[Top.scala 58:20]
  wire [15:0] n5_I_1; // @[Top.scala 58:20]
  wire [15:0] n5_I_2; // @[Top.scala 58:20]
  wire [15:0] n5_I_3; // @[Top.scala 58:20]
  wire [15:0] n5_I_4; // @[Top.scala 58:20]
  wire [15:0] n5_I_5; // @[Top.scala 58:20]
  wire [15:0] n5_I_6; // @[Top.scala 58:20]
  wire [15:0] n5_I_7; // @[Top.scala 58:20]
  wire [15:0] n5_I_8; // @[Top.scala 58:20]
  wire [15:0] n5_I_9; // @[Top.scala 58:20]
  wire [15:0] n5_I_10; // @[Top.scala 58:20]
  wire [15:0] n5_I_11; // @[Top.scala 58:20]
  wire [15:0] n5_I_12; // @[Top.scala 58:20]
  wire [15:0] n5_I_13; // @[Top.scala 58:20]
  wire [15:0] n5_I_14; // @[Top.scala 58:20]
  wire [15:0] n5_I_15; // @[Top.scala 58:20]
  wire [15:0] n5_O_0; // @[Top.scala 58:20]
  wire [15:0] n5_O_1; // @[Top.scala 58:20]
  wire [15:0] n5_O_2; // @[Top.scala 58:20]
  wire [15:0] n5_O_3; // @[Top.scala 58:20]
  wire [15:0] n5_O_4; // @[Top.scala 58:20]
  wire [15:0] n5_O_5; // @[Top.scala 58:20]
  wire [15:0] n5_O_6; // @[Top.scala 58:20]
  wire [15:0] n5_O_7; // @[Top.scala 58:20]
  wire [15:0] n5_O_8; // @[Top.scala 58:20]
  wire [15:0] n5_O_9; // @[Top.scala 58:20]
  wire [15:0] n5_O_10; // @[Top.scala 58:20]
  wire [15:0] n5_O_11; // @[Top.scala 58:20]
  wire [15:0] n5_O_12; // @[Top.scala 58:20]
  wire [15:0] n5_O_13; // @[Top.scala 58:20]
  wire [15:0] n5_O_14; // @[Top.scala 58:20]
  wire [15:0] n5_O_15; // @[Top.scala 58:20]
  wire  n6_clock; // @[Top.scala 61:20]
  wire  n6_reset; // @[Top.scala 61:20]
  wire  n6_valid_up; // @[Top.scala 61:20]
  wire  n6_valid_down; // @[Top.scala 61:20]
  wire [15:0] n6_I_0; // @[Top.scala 61:20]
  wire [15:0] n6_I_1; // @[Top.scala 61:20]
  wire [15:0] n6_I_2; // @[Top.scala 61:20]
  wire [15:0] n6_I_3; // @[Top.scala 61:20]
  wire [15:0] n6_I_4; // @[Top.scala 61:20]
  wire [15:0] n6_I_5; // @[Top.scala 61:20]
  wire [15:0] n6_I_6; // @[Top.scala 61:20]
  wire [15:0] n6_I_7; // @[Top.scala 61:20]
  wire [15:0] n6_I_8; // @[Top.scala 61:20]
  wire [15:0] n6_I_9; // @[Top.scala 61:20]
  wire [15:0] n6_I_10; // @[Top.scala 61:20]
  wire [15:0] n6_I_11; // @[Top.scala 61:20]
  wire [15:0] n6_I_12; // @[Top.scala 61:20]
  wire [15:0] n6_I_13; // @[Top.scala 61:20]
  wire [15:0] n6_I_14; // @[Top.scala 61:20]
  wire [15:0] n6_I_15; // @[Top.scala 61:20]
  wire [15:0] n6_O_0; // @[Top.scala 61:20]
  wire [15:0] n6_O_1; // @[Top.scala 61:20]
  wire [15:0] n6_O_2; // @[Top.scala 61:20]
  wire [15:0] n6_O_3; // @[Top.scala 61:20]
  wire [15:0] n6_O_4; // @[Top.scala 61:20]
  wire [15:0] n6_O_5; // @[Top.scala 61:20]
  wire [15:0] n6_O_6; // @[Top.scala 61:20]
  wire [15:0] n6_O_7; // @[Top.scala 61:20]
  wire [15:0] n6_O_8; // @[Top.scala 61:20]
  wire [15:0] n6_O_9; // @[Top.scala 61:20]
  wire [15:0] n6_O_10; // @[Top.scala 61:20]
  wire [15:0] n6_O_11; // @[Top.scala 61:20]
  wire [15:0] n6_O_12; // @[Top.scala 61:20]
  wire [15:0] n6_O_13; // @[Top.scala 61:20]
  wire [15:0] n6_O_14; // @[Top.scala 61:20]
  wire [15:0] n6_O_15; // @[Top.scala 61:20]
  wire  n7_valid_up; // @[Top.scala 64:20]
  wire  n7_valid_down; // @[Top.scala 64:20]
  wire [15:0] n7_I0_0; // @[Top.scala 64:20]
  wire [15:0] n7_I0_1; // @[Top.scala 64:20]
  wire [15:0] n7_I0_2; // @[Top.scala 64:20]
  wire [15:0] n7_I0_3; // @[Top.scala 64:20]
  wire [15:0] n7_I0_4; // @[Top.scala 64:20]
  wire [15:0] n7_I0_5; // @[Top.scala 64:20]
  wire [15:0] n7_I0_6; // @[Top.scala 64:20]
  wire [15:0] n7_I0_7; // @[Top.scala 64:20]
  wire [15:0] n7_I0_8; // @[Top.scala 64:20]
  wire [15:0] n7_I0_9; // @[Top.scala 64:20]
  wire [15:0] n7_I0_10; // @[Top.scala 64:20]
  wire [15:0] n7_I0_11; // @[Top.scala 64:20]
  wire [15:0] n7_I0_12; // @[Top.scala 64:20]
  wire [15:0] n7_I0_13; // @[Top.scala 64:20]
  wire [15:0] n7_I0_14; // @[Top.scala 64:20]
  wire [15:0] n7_I0_15; // @[Top.scala 64:20]
  wire [15:0] n7_I1_0; // @[Top.scala 64:20]
  wire [15:0] n7_I1_1; // @[Top.scala 64:20]
  wire [15:0] n7_I1_2; // @[Top.scala 64:20]
  wire [15:0] n7_I1_3; // @[Top.scala 64:20]
  wire [15:0] n7_I1_4; // @[Top.scala 64:20]
  wire [15:0] n7_I1_5; // @[Top.scala 64:20]
  wire [15:0] n7_I1_6; // @[Top.scala 64:20]
  wire [15:0] n7_I1_7; // @[Top.scala 64:20]
  wire [15:0] n7_I1_8; // @[Top.scala 64:20]
  wire [15:0] n7_I1_9; // @[Top.scala 64:20]
  wire [15:0] n7_I1_10; // @[Top.scala 64:20]
  wire [15:0] n7_I1_11; // @[Top.scala 64:20]
  wire [15:0] n7_I1_12; // @[Top.scala 64:20]
  wire [15:0] n7_I1_13; // @[Top.scala 64:20]
  wire [15:0] n7_I1_14; // @[Top.scala 64:20]
  wire [15:0] n7_I1_15; // @[Top.scala 64:20]
  wire [15:0] n7_O_0_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_0_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_1_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_1_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_2_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_2_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_3_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_3_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_4_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_4_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_5_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_5_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_6_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_6_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_7_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_7_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_8_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_8_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_9_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_9_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_10_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_10_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_11_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_11_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_12_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_12_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_13_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_13_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_14_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_14_1; // @[Top.scala 64:20]
  wire [15:0] n7_O_15_0; // @[Top.scala 64:20]
  wire [15:0] n7_O_15_1; // @[Top.scala 64:20]
  wire  n14_clock; // @[Top.scala 68:21]
  wire  n14_reset; // @[Top.scala 68:21]
  wire  n14_valid_up; // @[Top.scala 68:21]
  wire  n14_valid_down; // @[Top.scala 68:21]
  wire [15:0] n14_I_0; // @[Top.scala 68:21]
  wire [15:0] n14_I_1; // @[Top.scala 68:21]
  wire [15:0] n14_I_2; // @[Top.scala 68:21]
  wire [15:0] n14_I_3; // @[Top.scala 68:21]
  wire [15:0] n14_I_4; // @[Top.scala 68:21]
  wire [15:0] n14_I_5; // @[Top.scala 68:21]
  wire [15:0] n14_I_6; // @[Top.scala 68:21]
  wire [15:0] n14_I_7; // @[Top.scala 68:21]
  wire [15:0] n14_I_8; // @[Top.scala 68:21]
  wire [15:0] n14_I_9; // @[Top.scala 68:21]
  wire [15:0] n14_I_10; // @[Top.scala 68:21]
  wire [15:0] n14_I_11; // @[Top.scala 68:21]
  wire [15:0] n14_I_12; // @[Top.scala 68:21]
  wire [15:0] n14_I_13; // @[Top.scala 68:21]
  wire [15:0] n14_I_14; // @[Top.scala 68:21]
  wire [15:0] n14_I_15; // @[Top.scala 68:21]
  wire [15:0] n14_O_0; // @[Top.scala 68:21]
  wire [15:0] n14_O_1; // @[Top.scala 68:21]
  wire [15:0] n14_O_2; // @[Top.scala 68:21]
  wire [15:0] n14_O_3; // @[Top.scala 68:21]
  wire [15:0] n14_O_4; // @[Top.scala 68:21]
  wire [15:0] n14_O_5; // @[Top.scala 68:21]
  wire [15:0] n14_O_6; // @[Top.scala 68:21]
  wire [15:0] n14_O_7; // @[Top.scala 68:21]
  wire [15:0] n14_O_8; // @[Top.scala 68:21]
  wire [15:0] n14_O_9; // @[Top.scala 68:21]
  wire [15:0] n14_O_10; // @[Top.scala 68:21]
  wire [15:0] n14_O_11; // @[Top.scala 68:21]
  wire [15:0] n14_O_12; // @[Top.scala 68:21]
  wire [15:0] n14_O_13; // @[Top.scala 68:21]
  wire [15:0] n14_O_14; // @[Top.scala 68:21]
  wire [15:0] n14_O_15; // @[Top.scala 68:21]
  wire  n15_valid_up; // @[Top.scala 71:21]
  wire  n15_valid_down; // @[Top.scala 71:21]
  wire [15:0] n15_I0_0_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_0_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_1_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_1_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_2_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_2_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_3_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_3_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_4_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_4_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_5_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_5_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_6_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_6_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_7_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_7_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_8_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_8_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_9_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_9_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_10_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_10_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_11_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_11_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_12_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_12_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_13_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_13_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_14_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_14_1; // @[Top.scala 71:21]
  wire [15:0] n15_I0_15_0; // @[Top.scala 71:21]
  wire [15:0] n15_I0_15_1; // @[Top.scala 71:21]
  wire [15:0] n15_I1_0; // @[Top.scala 71:21]
  wire [15:0] n15_I1_1; // @[Top.scala 71:21]
  wire [15:0] n15_I1_2; // @[Top.scala 71:21]
  wire [15:0] n15_I1_3; // @[Top.scala 71:21]
  wire [15:0] n15_I1_4; // @[Top.scala 71:21]
  wire [15:0] n15_I1_5; // @[Top.scala 71:21]
  wire [15:0] n15_I1_6; // @[Top.scala 71:21]
  wire [15:0] n15_I1_7; // @[Top.scala 71:21]
  wire [15:0] n15_I1_8; // @[Top.scala 71:21]
  wire [15:0] n15_I1_9; // @[Top.scala 71:21]
  wire [15:0] n15_I1_10; // @[Top.scala 71:21]
  wire [15:0] n15_I1_11; // @[Top.scala 71:21]
  wire [15:0] n15_I1_12; // @[Top.scala 71:21]
  wire [15:0] n15_I1_13; // @[Top.scala 71:21]
  wire [15:0] n15_I1_14; // @[Top.scala 71:21]
  wire [15:0] n15_I1_15; // @[Top.scala 71:21]
  wire [15:0] n15_O_0_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_0_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_0_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_1_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_1_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_1_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_2_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_2_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_2_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_3_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_3_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_3_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_4_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_4_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_4_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_5_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_5_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_5_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_6_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_6_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_6_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_7_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_7_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_7_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_8_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_8_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_8_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_9_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_9_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_9_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_10_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_10_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_10_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_11_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_11_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_11_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_12_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_12_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_12_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_13_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_13_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_13_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_14_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_14_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_14_2; // @[Top.scala 71:21]
  wire [15:0] n15_O_15_0; // @[Top.scala 71:21]
  wire [15:0] n15_O_15_1; // @[Top.scala 71:21]
  wire [15:0] n15_O_15_2; // @[Top.scala 71:21]
  wire  n24_valid_up; // @[Top.scala 75:21]
  wire  n24_valid_down; // @[Top.scala 75:21]
  wire [15:0] n24_I_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_1_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_1_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_1_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_2_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_2_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_2_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_3_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_3_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_3_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_4_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_4_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_4_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_5_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_5_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_5_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_6_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_6_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_6_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_7_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_7_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_7_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_8_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_8_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_8_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_9_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_9_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_9_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_10_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_10_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_10_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_11_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_11_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_11_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_12_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_12_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_12_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_13_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_13_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_13_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_14_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_14_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_14_2; // @[Top.scala 75:21]
  wire [15:0] n24_I_15_0; // @[Top.scala 75:21]
  wire [15:0] n24_I_15_1; // @[Top.scala 75:21]
  wire [15:0] n24_I_15_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_0_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_0_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_0_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_1_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_1_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_1_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_2_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_2_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_2_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_3_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_3_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_3_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_4_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_4_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_4_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_5_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_5_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_5_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_6_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_6_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_6_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_7_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_7_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_7_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_8_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_8_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_8_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_9_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_9_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_9_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_10_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_10_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_10_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_11_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_11_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_11_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_12_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_12_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_12_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_13_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_13_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_13_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_14_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_14_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_14_0_2; // @[Top.scala 75:21]
  wire [15:0] n24_O_15_0_0; // @[Top.scala 75:21]
  wire [15:0] n24_O_15_0_1; // @[Top.scala 75:21]
  wire [15:0] n24_O_15_0_2; // @[Top.scala 75:21]
  wire  n31_valid_up; // @[Top.scala 78:21]
  wire  n31_valid_down; // @[Top.scala 78:21]
  wire [15:0] n31_I_0_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_0_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_0_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_1_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_1_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_1_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_2_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_2_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_2_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_3_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_3_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_3_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_4_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_4_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_4_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_5_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_5_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_5_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_6_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_6_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_6_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_7_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_7_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_7_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_8_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_8_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_8_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_9_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_9_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_9_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_10_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_10_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_10_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_11_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_11_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_11_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_12_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_12_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_12_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_13_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_13_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_13_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_14_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_14_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_14_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_I_15_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_I_15_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_I_15_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_0_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_0_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_0_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_1_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_1_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_1_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_2_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_2_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_2_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_3_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_3_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_3_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_4_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_4_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_4_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_5_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_5_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_5_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_6_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_6_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_6_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_7_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_7_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_7_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_8_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_8_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_8_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_9_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_9_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_9_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_10_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_10_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_10_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_11_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_11_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_11_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_12_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_12_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_12_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_13_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_13_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_13_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_14_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_14_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_14_2; // @[Top.scala 78:21]
  wire [15:0] n31_O_15_0; // @[Top.scala 78:21]
  wire [15:0] n31_O_15_1; // @[Top.scala 78:21]
  wire [15:0] n31_O_15_2; // @[Top.scala 78:21]
  wire  n32_clock; // @[Top.scala 81:21]
  wire  n32_reset; // @[Top.scala 81:21]
  wire  n32_valid_up; // @[Top.scala 81:21]
  wire  n32_valid_down; // @[Top.scala 81:21]
  wire [15:0] n32_I_0; // @[Top.scala 81:21]
  wire [15:0] n32_I_1; // @[Top.scala 81:21]
  wire [15:0] n32_I_2; // @[Top.scala 81:21]
  wire [15:0] n32_I_3; // @[Top.scala 81:21]
  wire [15:0] n32_I_4; // @[Top.scala 81:21]
  wire [15:0] n32_I_5; // @[Top.scala 81:21]
  wire [15:0] n32_I_6; // @[Top.scala 81:21]
  wire [15:0] n32_I_7; // @[Top.scala 81:21]
  wire [15:0] n32_I_8; // @[Top.scala 81:21]
  wire [15:0] n32_I_9; // @[Top.scala 81:21]
  wire [15:0] n32_I_10; // @[Top.scala 81:21]
  wire [15:0] n32_I_11; // @[Top.scala 81:21]
  wire [15:0] n32_I_12; // @[Top.scala 81:21]
  wire [15:0] n32_I_13; // @[Top.scala 81:21]
  wire [15:0] n32_I_14; // @[Top.scala 81:21]
  wire [15:0] n32_I_15; // @[Top.scala 81:21]
  wire [15:0] n32_O_0; // @[Top.scala 81:21]
  wire [15:0] n32_O_1; // @[Top.scala 81:21]
  wire [15:0] n32_O_2; // @[Top.scala 81:21]
  wire [15:0] n32_O_3; // @[Top.scala 81:21]
  wire [15:0] n32_O_4; // @[Top.scala 81:21]
  wire [15:0] n32_O_5; // @[Top.scala 81:21]
  wire [15:0] n32_O_6; // @[Top.scala 81:21]
  wire [15:0] n32_O_7; // @[Top.scala 81:21]
  wire [15:0] n32_O_8; // @[Top.scala 81:21]
  wire [15:0] n32_O_9; // @[Top.scala 81:21]
  wire [15:0] n32_O_10; // @[Top.scala 81:21]
  wire [15:0] n32_O_11; // @[Top.scala 81:21]
  wire [15:0] n32_O_12; // @[Top.scala 81:21]
  wire [15:0] n32_O_13; // @[Top.scala 81:21]
  wire [15:0] n32_O_14; // @[Top.scala 81:21]
  wire [15:0] n32_O_15; // @[Top.scala 81:21]
  wire  n33_clock; // @[Top.scala 84:21]
  wire  n33_reset; // @[Top.scala 84:21]
  wire  n33_valid_up; // @[Top.scala 84:21]
  wire  n33_valid_down; // @[Top.scala 84:21]
  wire [15:0] n33_I_0; // @[Top.scala 84:21]
  wire [15:0] n33_I_1; // @[Top.scala 84:21]
  wire [15:0] n33_I_2; // @[Top.scala 84:21]
  wire [15:0] n33_I_3; // @[Top.scala 84:21]
  wire [15:0] n33_I_4; // @[Top.scala 84:21]
  wire [15:0] n33_I_5; // @[Top.scala 84:21]
  wire [15:0] n33_I_6; // @[Top.scala 84:21]
  wire [15:0] n33_I_7; // @[Top.scala 84:21]
  wire [15:0] n33_I_8; // @[Top.scala 84:21]
  wire [15:0] n33_I_9; // @[Top.scala 84:21]
  wire [15:0] n33_I_10; // @[Top.scala 84:21]
  wire [15:0] n33_I_11; // @[Top.scala 84:21]
  wire [15:0] n33_I_12; // @[Top.scala 84:21]
  wire [15:0] n33_I_13; // @[Top.scala 84:21]
  wire [15:0] n33_I_14; // @[Top.scala 84:21]
  wire [15:0] n33_I_15; // @[Top.scala 84:21]
  wire [15:0] n33_O_0; // @[Top.scala 84:21]
  wire [15:0] n33_O_1; // @[Top.scala 84:21]
  wire [15:0] n33_O_2; // @[Top.scala 84:21]
  wire [15:0] n33_O_3; // @[Top.scala 84:21]
  wire [15:0] n33_O_4; // @[Top.scala 84:21]
  wire [15:0] n33_O_5; // @[Top.scala 84:21]
  wire [15:0] n33_O_6; // @[Top.scala 84:21]
  wire [15:0] n33_O_7; // @[Top.scala 84:21]
  wire [15:0] n33_O_8; // @[Top.scala 84:21]
  wire [15:0] n33_O_9; // @[Top.scala 84:21]
  wire [15:0] n33_O_10; // @[Top.scala 84:21]
  wire [15:0] n33_O_11; // @[Top.scala 84:21]
  wire [15:0] n33_O_12; // @[Top.scala 84:21]
  wire [15:0] n33_O_13; // @[Top.scala 84:21]
  wire [15:0] n33_O_14; // @[Top.scala 84:21]
  wire [15:0] n33_O_15; // @[Top.scala 84:21]
  wire  n34_clock; // @[Top.scala 87:21]
  wire  n34_reset; // @[Top.scala 87:21]
  wire  n34_valid_up; // @[Top.scala 87:21]
  wire  n34_valid_down; // @[Top.scala 87:21]
  wire [15:0] n34_I_0; // @[Top.scala 87:21]
  wire [15:0] n34_I_1; // @[Top.scala 87:21]
  wire [15:0] n34_I_2; // @[Top.scala 87:21]
  wire [15:0] n34_I_3; // @[Top.scala 87:21]
  wire [15:0] n34_I_4; // @[Top.scala 87:21]
  wire [15:0] n34_I_5; // @[Top.scala 87:21]
  wire [15:0] n34_I_6; // @[Top.scala 87:21]
  wire [15:0] n34_I_7; // @[Top.scala 87:21]
  wire [15:0] n34_I_8; // @[Top.scala 87:21]
  wire [15:0] n34_I_9; // @[Top.scala 87:21]
  wire [15:0] n34_I_10; // @[Top.scala 87:21]
  wire [15:0] n34_I_11; // @[Top.scala 87:21]
  wire [15:0] n34_I_12; // @[Top.scala 87:21]
  wire [15:0] n34_I_13; // @[Top.scala 87:21]
  wire [15:0] n34_I_14; // @[Top.scala 87:21]
  wire [15:0] n34_I_15; // @[Top.scala 87:21]
  wire [15:0] n34_O_0; // @[Top.scala 87:21]
  wire [15:0] n34_O_1; // @[Top.scala 87:21]
  wire [15:0] n34_O_2; // @[Top.scala 87:21]
  wire [15:0] n34_O_3; // @[Top.scala 87:21]
  wire [15:0] n34_O_4; // @[Top.scala 87:21]
  wire [15:0] n34_O_5; // @[Top.scala 87:21]
  wire [15:0] n34_O_6; // @[Top.scala 87:21]
  wire [15:0] n34_O_7; // @[Top.scala 87:21]
  wire [15:0] n34_O_8; // @[Top.scala 87:21]
  wire [15:0] n34_O_9; // @[Top.scala 87:21]
  wire [15:0] n34_O_10; // @[Top.scala 87:21]
  wire [15:0] n34_O_11; // @[Top.scala 87:21]
  wire [15:0] n34_O_12; // @[Top.scala 87:21]
  wire [15:0] n34_O_13; // @[Top.scala 87:21]
  wire [15:0] n34_O_14; // @[Top.scala 87:21]
  wire [15:0] n34_O_15; // @[Top.scala 87:21]
  wire  n35_valid_up; // @[Top.scala 90:21]
  wire  n35_valid_down; // @[Top.scala 90:21]
  wire [15:0] n35_I0_0; // @[Top.scala 90:21]
  wire [15:0] n35_I0_1; // @[Top.scala 90:21]
  wire [15:0] n35_I0_2; // @[Top.scala 90:21]
  wire [15:0] n35_I0_3; // @[Top.scala 90:21]
  wire [15:0] n35_I0_4; // @[Top.scala 90:21]
  wire [15:0] n35_I0_5; // @[Top.scala 90:21]
  wire [15:0] n35_I0_6; // @[Top.scala 90:21]
  wire [15:0] n35_I0_7; // @[Top.scala 90:21]
  wire [15:0] n35_I0_8; // @[Top.scala 90:21]
  wire [15:0] n35_I0_9; // @[Top.scala 90:21]
  wire [15:0] n35_I0_10; // @[Top.scala 90:21]
  wire [15:0] n35_I0_11; // @[Top.scala 90:21]
  wire [15:0] n35_I0_12; // @[Top.scala 90:21]
  wire [15:0] n35_I0_13; // @[Top.scala 90:21]
  wire [15:0] n35_I0_14; // @[Top.scala 90:21]
  wire [15:0] n35_I0_15; // @[Top.scala 90:21]
  wire [15:0] n35_I1_0; // @[Top.scala 90:21]
  wire [15:0] n35_I1_1; // @[Top.scala 90:21]
  wire [15:0] n35_I1_2; // @[Top.scala 90:21]
  wire [15:0] n35_I1_3; // @[Top.scala 90:21]
  wire [15:0] n35_I1_4; // @[Top.scala 90:21]
  wire [15:0] n35_I1_5; // @[Top.scala 90:21]
  wire [15:0] n35_I1_6; // @[Top.scala 90:21]
  wire [15:0] n35_I1_7; // @[Top.scala 90:21]
  wire [15:0] n35_I1_8; // @[Top.scala 90:21]
  wire [15:0] n35_I1_9; // @[Top.scala 90:21]
  wire [15:0] n35_I1_10; // @[Top.scala 90:21]
  wire [15:0] n35_I1_11; // @[Top.scala 90:21]
  wire [15:0] n35_I1_12; // @[Top.scala 90:21]
  wire [15:0] n35_I1_13; // @[Top.scala 90:21]
  wire [15:0] n35_I1_14; // @[Top.scala 90:21]
  wire [15:0] n35_I1_15; // @[Top.scala 90:21]
  wire [15:0] n35_O_0_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_0_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_1_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_1_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_2_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_2_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_3_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_3_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_4_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_4_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_5_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_5_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_6_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_6_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_7_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_7_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_8_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_8_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_9_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_9_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_10_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_10_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_11_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_11_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_12_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_12_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_13_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_13_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_14_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_14_1; // @[Top.scala 90:21]
  wire [15:0] n35_O_15_0; // @[Top.scala 90:21]
  wire [15:0] n35_O_15_1; // @[Top.scala 90:21]
  wire  n42_clock; // @[Top.scala 94:21]
  wire  n42_reset; // @[Top.scala 94:21]
  wire  n42_valid_up; // @[Top.scala 94:21]
  wire  n42_valid_down; // @[Top.scala 94:21]
  wire [15:0] n42_I_0; // @[Top.scala 94:21]
  wire [15:0] n42_I_1; // @[Top.scala 94:21]
  wire [15:0] n42_I_2; // @[Top.scala 94:21]
  wire [15:0] n42_I_3; // @[Top.scala 94:21]
  wire [15:0] n42_I_4; // @[Top.scala 94:21]
  wire [15:0] n42_I_5; // @[Top.scala 94:21]
  wire [15:0] n42_I_6; // @[Top.scala 94:21]
  wire [15:0] n42_I_7; // @[Top.scala 94:21]
  wire [15:0] n42_I_8; // @[Top.scala 94:21]
  wire [15:0] n42_I_9; // @[Top.scala 94:21]
  wire [15:0] n42_I_10; // @[Top.scala 94:21]
  wire [15:0] n42_I_11; // @[Top.scala 94:21]
  wire [15:0] n42_I_12; // @[Top.scala 94:21]
  wire [15:0] n42_I_13; // @[Top.scala 94:21]
  wire [15:0] n42_I_14; // @[Top.scala 94:21]
  wire [15:0] n42_I_15; // @[Top.scala 94:21]
  wire [15:0] n42_O_0; // @[Top.scala 94:21]
  wire [15:0] n42_O_1; // @[Top.scala 94:21]
  wire [15:0] n42_O_2; // @[Top.scala 94:21]
  wire [15:0] n42_O_3; // @[Top.scala 94:21]
  wire [15:0] n42_O_4; // @[Top.scala 94:21]
  wire [15:0] n42_O_5; // @[Top.scala 94:21]
  wire [15:0] n42_O_6; // @[Top.scala 94:21]
  wire [15:0] n42_O_7; // @[Top.scala 94:21]
  wire [15:0] n42_O_8; // @[Top.scala 94:21]
  wire [15:0] n42_O_9; // @[Top.scala 94:21]
  wire [15:0] n42_O_10; // @[Top.scala 94:21]
  wire [15:0] n42_O_11; // @[Top.scala 94:21]
  wire [15:0] n42_O_12; // @[Top.scala 94:21]
  wire [15:0] n42_O_13; // @[Top.scala 94:21]
  wire [15:0] n42_O_14; // @[Top.scala 94:21]
  wire [15:0] n42_O_15; // @[Top.scala 94:21]
  wire  n43_valid_up; // @[Top.scala 97:21]
  wire  n43_valid_down; // @[Top.scala 97:21]
  wire [15:0] n43_I0_0_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_0_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_1_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_1_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_2_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_2_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_3_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_3_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_4_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_4_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_5_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_5_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_6_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_6_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_7_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_7_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_8_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_8_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_9_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_9_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_10_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_10_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_11_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_11_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_12_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_12_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_13_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_13_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_14_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_14_1; // @[Top.scala 97:21]
  wire [15:0] n43_I0_15_0; // @[Top.scala 97:21]
  wire [15:0] n43_I0_15_1; // @[Top.scala 97:21]
  wire [15:0] n43_I1_0; // @[Top.scala 97:21]
  wire [15:0] n43_I1_1; // @[Top.scala 97:21]
  wire [15:0] n43_I1_2; // @[Top.scala 97:21]
  wire [15:0] n43_I1_3; // @[Top.scala 97:21]
  wire [15:0] n43_I1_4; // @[Top.scala 97:21]
  wire [15:0] n43_I1_5; // @[Top.scala 97:21]
  wire [15:0] n43_I1_6; // @[Top.scala 97:21]
  wire [15:0] n43_I1_7; // @[Top.scala 97:21]
  wire [15:0] n43_I1_8; // @[Top.scala 97:21]
  wire [15:0] n43_I1_9; // @[Top.scala 97:21]
  wire [15:0] n43_I1_10; // @[Top.scala 97:21]
  wire [15:0] n43_I1_11; // @[Top.scala 97:21]
  wire [15:0] n43_I1_12; // @[Top.scala 97:21]
  wire [15:0] n43_I1_13; // @[Top.scala 97:21]
  wire [15:0] n43_I1_14; // @[Top.scala 97:21]
  wire [15:0] n43_I1_15; // @[Top.scala 97:21]
  wire [15:0] n43_O_0_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_0_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_0_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_1_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_1_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_1_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_2_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_2_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_2_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_3_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_3_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_3_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_4_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_4_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_4_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_5_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_5_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_5_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_6_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_6_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_6_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_7_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_7_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_7_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_8_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_8_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_8_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_9_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_9_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_9_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_10_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_10_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_10_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_11_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_11_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_11_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_12_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_12_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_12_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_13_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_13_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_13_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_14_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_14_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_14_2; // @[Top.scala 97:21]
  wire [15:0] n43_O_15_0; // @[Top.scala 97:21]
  wire [15:0] n43_O_15_1; // @[Top.scala 97:21]
  wire [15:0] n43_O_15_2; // @[Top.scala 97:21]
  wire  n52_valid_up; // @[Top.scala 101:21]
  wire  n52_valid_down; // @[Top.scala 101:21]
  wire [15:0] n52_I_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_1_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_1_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_1_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_2_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_2_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_2_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_3_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_3_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_3_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_4_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_4_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_4_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_5_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_5_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_5_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_6_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_6_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_6_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_7_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_7_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_7_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_8_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_8_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_8_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_9_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_9_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_9_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_10_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_10_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_10_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_11_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_11_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_11_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_12_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_12_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_12_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_13_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_13_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_13_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_14_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_14_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_14_2; // @[Top.scala 101:21]
  wire [15:0] n52_I_15_0; // @[Top.scala 101:21]
  wire [15:0] n52_I_15_1; // @[Top.scala 101:21]
  wire [15:0] n52_I_15_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_0_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_0_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_0_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_1_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_1_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_1_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_2_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_2_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_2_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_3_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_3_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_3_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_4_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_4_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_4_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_5_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_5_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_5_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_6_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_6_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_6_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_7_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_7_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_7_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_8_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_8_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_8_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_9_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_9_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_9_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_10_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_10_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_10_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_11_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_11_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_11_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_12_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_12_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_12_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_13_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_13_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_13_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_14_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_14_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_14_0_2; // @[Top.scala 101:21]
  wire [15:0] n52_O_15_0_0; // @[Top.scala 101:21]
  wire [15:0] n52_O_15_0_1; // @[Top.scala 101:21]
  wire [15:0] n52_O_15_0_2; // @[Top.scala 101:21]
  wire  n59_valid_up; // @[Top.scala 104:21]
  wire  n59_valid_down; // @[Top.scala 104:21]
  wire [15:0] n59_I_0_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_0_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_0_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_1_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_1_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_1_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_2_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_2_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_2_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_3_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_3_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_3_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_4_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_4_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_4_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_5_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_5_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_5_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_6_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_6_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_6_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_7_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_7_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_7_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_8_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_8_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_8_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_9_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_9_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_9_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_10_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_10_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_10_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_11_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_11_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_11_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_12_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_12_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_12_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_13_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_13_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_13_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_14_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_14_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_14_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_I_15_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_I_15_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_I_15_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_0_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_0_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_0_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_1_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_1_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_1_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_2_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_2_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_2_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_3_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_3_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_3_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_4_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_4_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_4_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_5_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_5_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_5_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_6_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_6_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_6_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_7_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_7_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_7_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_8_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_8_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_8_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_9_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_9_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_9_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_10_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_10_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_10_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_11_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_11_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_11_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_12_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_12_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_12_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_13_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_13_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_13_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_14_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_14_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_14_2; // @[Top.scala 104:21]
  wire [15:0] n59_O_15_0; // @[Top.scala 104:21]
  wire [15:0] n59_O_15_1; // @[Top.scala 104:21]
  wire [15:0] n59_O_15_2; // @[Top.scala 104:21]
  wire  n60_clock; // @[Top.scala 107:21]
  wire  n60_reset; // @[Top.scala 107:21]
  wire  n60_valid_up; // @[Top.scala 107:21]
  wire  n60_valid_down; // @[Top.scala 107:21]
  wire [15:0] n60_I_0_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_0_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_0_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_1_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_1_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_1_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_2_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_2_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_2_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_3_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_3_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_3_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_4_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_4_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_4_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_5_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_5_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_5_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_6_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_6_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_6_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_7_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_7_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_7_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_8_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_8_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_8_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_9_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_9_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_9_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_10_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_10_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_10_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_11_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_11_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_11_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_12_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_12_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_12_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_13_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_13_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_13_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_14_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_14_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_14_2; // @[Top.scala 107:21]
  wire [15:0] n60_I_15_0; // @[Top.scala 107:21]
  wire [15:0] n60_I_15_1; // @[Top.scala 107:21]
  wire [15:0] n60_I_15_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_0_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_0_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_0_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_1_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_1_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_1_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_2_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_2_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_2_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_3_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_3_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_3_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_4_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_4_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_4_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_5_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_5_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_5_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_6_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_6_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_6_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_7_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_7_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_7_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_8_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_8_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_8_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_9_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_9_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_9_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_10_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_10_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_10_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_11_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_11_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_11_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_12_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_12_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_12_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_13_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_13_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_13_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_14_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_14_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_14_2; // @[Top.scala 107:21]
  wire [15:0] n60_O_15_0; // @[Top.scala 107:21]
  wire [15:0] n60_O_15_1; // @[Top.scala 107:21]
  wire [15:0] n60_O_15_2; // @[Top.scala 107:21]
  wire  n61_valid_up; // @[Top.scala 110:21]
  wire  n61_valid_down; // @[Top.scala 110:21]
  wire [15:0] n61_I0_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_2_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_2_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_2_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_3_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_3_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_3_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_4_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_4_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_4_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_5_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_5_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_5_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_6_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_6_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_6_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_7_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_7_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_7_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_8_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_8_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_8_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_9_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_9_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_9_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_10_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_10_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_10_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_11_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_11_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_11_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_12_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_12_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_12_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_13_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_13_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_13_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_14_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_14_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_14_2; // @[Top.scala 110:21]
  wire [15:0] n61_I0_15_0; // @[Top.scala 110:21]
  wire [15:0] n61_I0_15_1; // @[Top.scala 110:21]
  wire [15:0] n61_I0_15_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_2_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_2_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_2_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_3_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_3_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_3_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_4_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_4_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_4_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_5_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_5_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_5_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_6_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_6_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_6_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_7_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_7_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_7_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_8_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_8_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_8_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_9_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_9_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_9_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_10_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_10_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_10_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_11_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_11_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_11_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_12_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_12_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_12_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_13_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_13_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_13_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_14_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_14_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_14_2; // @[Top.scala 110:21]
  wire [15:0] n61_I1_15_0; // @[Top.scala 110:21]
  wire [15:0] n61_I1_15_1; // @[Top.scala 110:21]
  wire [15:0] n61_I1_15_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_0_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_0_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_0_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_0_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_0_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_0_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_1_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_1_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_1_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_1_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_1_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_1_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_2_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_2_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_2_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_2_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_2_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_2_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_3_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_3_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_3_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_3_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_3_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_3_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_4_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_4_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_4_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_4_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_4_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_4_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_5_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_5_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_5_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_5_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_5_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_5_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_6_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_6_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_6_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_6_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_6_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_6_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_7_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_7_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_7_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_7_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_7_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_7_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_8_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_8_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_8_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_8_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_8_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_8_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_9_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_9_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_9_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_9_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_9_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_9_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_10_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_10_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_10_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_10_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_10_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_10_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_11_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_11_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_11_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_11_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_11_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_11_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_12_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_12_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_12_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_12_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_12_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_12_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_13_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_13_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_13_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_13_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_13_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_13_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_14_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_14_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_14_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_14_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_14_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_14_1_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_15_0_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_15_0_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_15_0_2; // @[Top.scala 110:21]
  wire [15:0] n61_O_15_1_0; // @[Top.scala 110:21]
  wire [15:0] n61_O_15_1_1; // @[Top.scala 110:21]
  wire [15:0] n61_O_15_1_2; // @[Top.scala 110:21]
  wire  n68_clock; // @[Top.scala 114:21]
  wire  n68_reset; // @[Top.scala 114:21]
  wire  n68_valid_up; // @[Top.scala 114:21]
  wire  n68_valid_down; // @[Top.scala 114:21]
  wire [15:0] n68_I_0; // @[Top.scala 114:21]
  wire [15:0] n68_I_1; // @[Top.scala 114:21]
  wire [15:0] n68_I_2; // @[Top.scala 114:21]
  wire [15:0] n68_I_3; // @[Top.scala 114:21]
  wire [15:0] n68_I_4; // @[Top.scala 114:21]
  wire [15:0] n68_I_5; // @[Top.scala 114:21]
  wire [15:0] n68_I_6; // @[Top.scala 114:21]
  wire [15:0] n68_I_7; // @[Top.scala 114:21]
  wire [15:0] n68_I_8; // @[Top.scala 114:21]
  wire [15:0] n68_I_9; // @[Top.scala 114:21]
  wire [15:0] n68_I_10; // @[Top.scala 114:21]
  wire [15:0] n68_I_11; // @[Top.scala 114:21]
  wire [15:0] n68_I_12; // @[Top.scala 114:21]
  wire [15:0] n68_I_13; // @[Top.scala 114:21]
  wire [15:0] n68_I_14; // @[Top.scala 114:21]
  wire [15:0] n68_I_15; // @[Top.scala 114:21]
  wire [15:0] n68_O_0; // @[Top.scala 114:21]
  wire [15:0] n68_O_1; // @[Top.scala 114:21]
  wire [15:0] n68_O_2; // @[Top.scala 114:21]
  wire [15:0] n68_O_3; // @[Top.scala 114:21]
  wire [15:0] n68_O_4; // @[Top.scala 114:21]
  wire [15:0] n68_O_5; // @[Top.scala 114:21]
  wire [15:0] n68_O_6; // @[Top.scala 114:21]
  wire [15:0] n68_O_7; // @[Top.scala 114:21]
  wire [15:0] n68_O_8; // @[Top.scala 114:21]
  wire [15:0] n68_O_9; // @[Top.scala 114:21]
  wire [15:0] n68_O_10; // @[Top.scala 114:21]
  wire [15:0] n68_O_11; // @[Top.scala 114:21]
  wire [15:0] n68_O_12; // @[Top.scala 114:21]
  wire [15:0] n68_O_13; // @[Top.scala 114:21]
  wire [15:0] n68_O_14; // @[Top.scala 114:21]
  wire [15:0] n68_O_15; // @[Top.scala 114:21]
  wire  n69_clock; // @[Top.scala 117:21]
  wire  n69_reset; // @[Top.scala 117:21]
  wire  n69_valid_up; // @[Top.scala 117:21]
  wire  n69_valid_down; // @[Top.scala 117:21]
  wire [15:0] n69_I_0; // @[Top.scala 117:21]
  wire [15:0] n69_I_1; // @[Top.scala 117:21]
  wire [15:0] n69_I_2; // @[Top.scala 117:21]
  wire [15:0] n69_I_3; // @[Top.scala 117:21]
  wire [15:0] n69_I_4; // @[Top.scala 117:21]
  wire [15:0] n69_I_5; // @[Top.scala 117:21]
  wire [15:0] n69_I_6; // @[Top.scala 117:21]
  wire [15:0] n69_I_7; // @[Top.scala 117:21]
  wire [15:0] n69_I_8; // @[Top.scala 117:21]
  wire [15:0] n69_I_9; // @[Top.scala 117:21]
  wire [15:0] n69_I_10; // @[Top.scala 117:21]
  wire [15:0] n69_I_11; // @[Top.scala 117:21]
  wire [15:0] n69_I_12; // @[Top.scala 117:21]
  wire [15:0] n69_I_13; // @[Top.scala 117:21]
  wire [15:0] n69_I_14; // @[Top.scala 117:21]
  wire [15:0] n69_I_15; // @[Top.scala 117:21]
  wire [15:0] n69_O_0; // @[Top.scala 117:21]
  wire [15:0] n69_O_1; // @[Top.scala 117:21]
  wire [15:0] n69_O_2; // @[Top.scala 117:21]
  wire [15:0] n69_O_3; // @[Top.scala 117:21]
  wire [15:0] n69_O_4; // @[Top.scala 117:21]
  wire [15:0] n69_O_5; // @[Top.scala 117:21]
  wire [15:0] n69_O_6; // @[Top.scala 117:21]
  wire [15:0] n69_O_7; // @[Top.scala 117:21]
  wire [15:0] n69_O_8; // @[Top.scala 117:21]
  wire [15:0] n69_O_9; // @[Top.scala 117:21]
  wire [15:0] n69_O_10; // @[Top.scala 117:21]
  wire [15:0] n69_O_11; // @[Top.scala 117:21]
  wire [15:0] n69_O_12; // @[Top.scala 117:21]
  wire [15:0] n69_O_13; // @[Top.scala 117:21]
  wire [15:0] n69_O_14; // @[Top.scala 117:21]
  wire [15:0] n69_O_15; // @[Top.scala 117:21]
  wire  n70_clock; // @[Top.scala 120:21]
  wire  n70_reset; // @[Top.scala 120:21]
  wire  n70_valid_up; // @[Top.scala 120:21]
  wire  n70_valid_down; // @[Top.scala 120:21]
  wire [15:0] n70_I_0; // @[Top.scala 120:21]
  wire [15:0] n70_I_1; // @[Top.scala 120:21]
  wire [15:0] n70_I_2; // @[Top.scala 120:21]
  wire [15:0] n70_I_3; // @[Top.scala 120:21]
  wire [15:0] n70_I_4; // @[Top.scala 120:21]
  wire [15:0] n70_I_5; // @[Top.scala 120:21]
  wire [15:0] n70_I_6; // @[Top.scala 120:21]
  wire [15:0] n70_I_7; // @[Top.scala 120:21]
  wire [15:0] n70_I_8; // @[Top.scala 120:21]
  wire [15:0] n70_I_9; // @[Top.scala 120:21]
  wire [15:0] n70_I_10; // @[Top.scala 120:21]
  wire [15:0] n70_I_11; // @[Top.scala 120:21]
  wire [15:0] n70_I_12; // @[Top.scala 120:21]
  wire [15:0] n70_I_13; // @[Top.scala 120:21]
  wire [15:0] n70_I_14; // @[Top.scala 120:21]
  wire [15:0] n70_I_15; // @[Top.scala 120:21]
  wire [15:0] n70_O_0; // @[Top.scala 120:21]
  wire [15:0] n70_O_1; // @[Top.scala 120:21]
  wire [15:0] n70_O_2; // @[Top.scala 120:21]
  wire [15:0] n70_O_3; // @[Top.scala 120:21]
  wire [15:0] n70_O_4; // @[Top.scala 120:21]
  wire [15:0] n70_O_5; // @[Top.scala 120:21]
  wire [15:0] n70_O_6; // @[Top.scala 120:21]
  wire [15:0] n70_O_7; // @[Top.scala 120:21]
  wire [15:0] n70_O_8; // @[Top.scala 120:21]
  wire [15:0] n70_O_9; // @[Top.scala 120:21]
  wire [15:0] n70_O_10; // @[Top.scala 120:21]
  wire [15:0] n70_O_11; // @[Top.scala 120:21]
  wire [15:0] n70_O_12; // @[Top.scala 120:21]
  wire [15:0] n70_O_13; // @[Top.scala 120:21]
  wire [15:0] n70_O_14; // @[Top.scala 120:21]
  wire [15:0] n70_O_15; // @[Top.scala 120:21]
  wire  n71_valid_up; // @[Top.scala 123:21]
  wire  n71_valid_down; // @[Top.scala 123:21]
  wire [15:0] n71_I0_0; // @[Top.scala 123:21]
  wire [15:0] n71_I0_1; // @[Top.scala 123:21]
  wire [15:0] n71_I0_2; // @[Top.scala 123:21]
  wire [15:0] n71_I0_3; // @[Top.scala 123:21]
  wire [15:0] n71_I0_4; // @[Top.scala 123:21]
  wire [15:0] n71_I0_5; // @[Top.scala 123:21]
  wire [15:0] n71_I0_6; // @[Top.scala 123:21]
  wire [15:0] n71_I0_7; // @[Top.scala 123:21]
  wire [15:0] n71_I0_8; // @[Top.scala 123:21]
  wire [15:0] n71_I0_9; // @[Top.scala 123:21]
  wire [15:0] n71_I0_10; // @[Top.scala 123:21]
  wire [15:0] n71_I0_11; // @[Top.scala 123:21]
  wire [15:0] n71_I0_12; // @[Top.scala 123:21]
  wire [15:0] n71_I0_13; // @[Top.scala 123:21]
  wire [15:0] n71_I0_14; // @[Top.scala 123:21]
  wire [15:0] n71_I0_15; // @[Top.scala 123:21]
  wire [15:0] n71_I1_0; // @[Top.scala 123:21]
  wire [15:0] n71_I1_1; // @[Top.scala 123:21]
  wire [15:0] n71_I1_2; // @[Top.scala 123:21]
  wire [15:0] n71_I1_3; // @[Top.scala 123:21]
  wire [15:0] n71_I1_4; // @[Top.scala 123:21]
  wire [15:0] n71_I1_5; // @[Top.scala 123:21]
  wire [15:0] n71_I1_6; // @[Top.scala 123:21]
  wire [15:0] n71_I1_7; // @[Top.scala 123:21]
  wire [15:0] n71_I1_8; // @[Top.scala 123:21]
  wire [15:0] n71_I1_9; // @[Top.scala 123:21]
  wire [15:0] n71_I1_10; // @[Top.scala 123:21]
  wire [15:0] n71_I1_11; // @[Top.scala 123:21]
  wire [15:0] n71_I1_12; // @[Top.scala 123:21]
  wire [15:0] n71_I1_13; // @[Top.scala 123:21]
  wire [15:0] n71_I1_14; // @[Top.scala 123:21]
  wire [15:0] n71_I1_15; // @[Top.scala 123:21]
  wire [15:0] n71_O_0_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_0_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_1_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_1_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_2_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_2_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_3_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_3_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_4_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_4_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_5_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_5_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_6_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_6_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_7_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_7_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_8_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_8_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_9_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_9_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_10_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_10_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_11_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_11_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_12_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_12_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_13_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_13_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_14_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_14_1; // @[Top.scala 123:21]
  wire [15:0] n71_O_15_0; // @[Top.scala 123:21]
  wire [15:0] n71_O_15_1; // @[Top.scala 123:21]
  wire  n78_clock; // @[Top.scala 127:21]
  wire  n78_reset; // @[Top.scala 127:21]
  wire  n78_valid_up; // @[Top.scala 127:21]
  wire  n78_valid_down; // @[Top.scala 127:21]
  wire [15:0] n78_I_0; // @[Top.scala 127:21]
  wire [15:0] n78_I_1; // @[Top.scala 127:21]
  wire [15:0] n78_I_2; // @[Top.scala 127:21]
  wire [15:0] n78_I_3; // @[Top.scala 127:21]
  wire [15:0] n78_I_4; // @[Top.scala 127:21]
  wire [15:0] n78_I_5; // @[Top.scala 127:21]
  wire [15:0] n78_I_6; // @[Top.scala 127:21]
  wire [15:0] n78_I_7; // @[Top.scala 127:21]
  wire [15:0] n78_I_8; // @[Top.scala 127:21]
  wire [15:0] n78_I_9; // @[Top.scala 127:21]
  wire [15:0] n78_I_10; // @[Top.scala 127:21]
  wire [15:0] n78_I_11; // @[Top.scala 127:21]
  wire [15:0] n78_I_12; // @[Top.scala 127:21]
  wire [15:0] n78_I_13; // @[Top.scala 127:21]
  wire [15:0] n78_I_14; // @[Top.scala 127:21]
  wire [15:0] n78_I_15; // @[Top.scala 127:21]
  wire [15:0] n78_O_0; // @[Top.scala 127:21]
  wire [15:0] n78_O_1; // @[Top.scala 127:21]
  wire [15:0] n78_O_2; // @[Top.scala 127:21]
  wire [15:0] n78_O_3; // @[Top.scala 127:21]
  wire [15:0] n78_O_4; // @[Top.scala 127:21]
  wire [15:0] n78_O_5; // @[Top.scala 127:21]
  wire [15:0] n78_O_6; // @[Top.scala 127:21]
  wire [15:0] n78_O_7; // @[Top.scala 127:21]
  wire [15:0] n78_O_8; // @[Top.scala 127:21]
  wire [15:0] n78_O_9; // @[Top.scala 127:21]
  wire [15:0] n78_O_10; // @[Top.scala 127:21]
  wire [15:0] n78_O_11; // @[Top.scala 127:21]
  wire [15:0] n78_O_12; // @[Top.scala 127:21]
  wire [15:0] n78_O_13; // @[Top.scala 127:21]
  wire [15:0] n78_O_14; // @[Top.scala 127:21]
  wire [15:0] n78_O_15; // @[Top.scala 127:21]
  wire  n79_valid_up; // @[Top.scala 130:21]
  wire  n79_valid_down; // @[Top.scala 130:21]
  wire [15:0] n79_I0_0_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_0_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_1_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_1_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_2_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_2_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_3_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_3_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_4_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_4_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_5_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_5_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_6_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_6_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_7_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_7_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_8_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_8_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_9_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_9_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_10_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_10_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_11_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_11_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_12_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_12_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_13_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_13_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_14_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_14_1; // @[Top.scala 130:21]
  wire [15:0] n79_I0_15_0; // @[Top.scala 130:21]
  wire [15:0] n79_I0_15_1; // @[Top.scala 130:21]
  wire [15:0] n79_I1_0; // @[Top.scala 130:21]
  wire [15:0] n79_I1_1; // @[Top.scala 130:21]
  wire [15:0] n79_I1_2; // @[Top.scala 130:21]
  wire [15:0] n79_I1_3; // @[Top.scala 130:21]
  wire [15:0] n79_I1_4; // @[Top.scala 130:21]
  wire [15:0] n79_I1_5; // @[Top.scala 130:21]
  wire [15:0] n79_I1_6; // @[Top.scala 130:21]
  wire [15:0] n79_I1_7; // @[Top.scala 130:21]
  wire [15:0] n79_I1_8; // @[Top.scala 130:21]
  wire [15:0] n79_I1_9; // @[Top.scala 130:21]
  wire [15:0] n79_I1_10; // @[Top.scala 130:21]
  wire [15:0] n79_I1_11; // @[Top.scala 130:21]
  wire [15:0] n79_I1_12; // @[Top.scala 130:21]
  wire [15:0] n79_I1_13; // @[Top.scala 130:21]
  wire [15:0] n79_I1_14; // @[Top.scala 130:21]
  wire [15:0] n79_I1_15; // @[Top.scala 130:21]
  wire [15:0] n79_O_0_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_0_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_0_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_1_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_1_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_1_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_2_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_2_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_2_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_3_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_3_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_3_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_4_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_4_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_4_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_5_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_5_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_5_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_6_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_6_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_6_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_7_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_7_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_7_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_8_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_8_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_8_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_9_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_9_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_9_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_10_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_10_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_10_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_11_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_11_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_11_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_12_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_12_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_12_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_13_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_13_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_13_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_14_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_14_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_14_2; // @[Top.scala 130:21]
  wire [15:0] n79_O_15_0; // @[Top.scala 130:21]
  wire [15:0] n79_O_15_1; // @[Top.scala 130:21]
  wire [15:0] n79_O_15_2; // @[Top.scala 130:21]
  wire  n88_valid_up; // @[Top.scala 134:21]
  wire  n88_valid_down; // @[Top.scala 134:21]
  wire [15:0] n88_I_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_1_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_1_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_1_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_2_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_2_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_2_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_3_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_3_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_3_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_4_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_4_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_4_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_5_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_5_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_5_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_6_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_6_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_6_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_7_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_7_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_7_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_8_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_8_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_8_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_9_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_9_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_9_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_10_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_10_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_10_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_11_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_11_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_11_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_12_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_12_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_12_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_13_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_13_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_13_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_14_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_14_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_14_2; // @[Top.scala 134:21]
  wire [15:0] n88_I_15_0; // @[Top.scala 134:21]
  wire [15:0] n88_I_15_1; // @[Top.scala 134:21]
  wire [15:0] n88_I_15_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_0_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_0_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_0_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_1_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_1_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_1_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_2_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_2_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_2_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_3_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_3_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_3_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_4_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_4_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_4_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_5_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_5_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_5_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_6_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_6_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_6_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_7_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_7_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_7_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_8_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_8_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_8_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_9_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_9_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_9_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_10_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_10_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_10_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_11_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_11_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_11_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_12_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_12_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_12_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_13_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_13_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_13_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_14_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_14_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_14_0_2; // @[Top.scala 134:21]
  wire [15:0] n88_O_15_0_0; // @[Top.scala 134:21]
  wire [15:0] n88_O_15_0_1; // @[Top.scala 134:21]
  wire [15:0] n88_O_15_0_2; // @[Top.scala 134:21]
  wire  n95_valid_up; // @[Top.scala 137:21]
  wire  n95_valid_down; // @[Top.scala 137:21]
  wire [15:0] n95_I_0_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_0_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_0_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_1_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_1_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_1_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_2_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_2_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_2_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_3_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_3_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_3_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_4_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_4_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_4_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_5_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_5_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_5_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_6_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_6_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_6_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_7_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_7_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_7_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_8_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_8_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_8_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_9_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_9_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_9_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_10_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_10_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_10_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_11_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_11_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_11_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_12_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_12_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_12_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_13_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_13_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_13_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_14_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_14_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_14_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_I_15_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_I_15_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_I_15_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_0_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_0_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_0_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_1_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_1_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_1_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_2_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_2_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_2_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_3_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_3_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_3_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_4_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_4_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_4_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_5_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_5_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_5_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_6_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_6_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_6_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_7_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_7_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_7_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_8_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_8_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_8_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_9_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_9_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_9_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_10_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_10_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_10_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_11_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_11_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_11_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_12_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_12_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_12_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_13_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_13_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_13_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_14_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_14_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_14_2; // @[Top.scala 137:21]
  wire [15:0] n95_O_15_0; // @[Top.scala 137:21]
  wire [15:0] n95_O_15_1; // @[Top.scala 137:21]
  wire [15:0] n95_O_15_2; // @[Top.scala 137:21]
  wire  n96_clock; // @[Top.scala 140:21]
  wire  n96_reset; // @[Top.scala 140:21]
  wire  n96_valid_up; // @[Top.scala 140:21]
  wire  n96_valid_down; // @[Top.scala 140:21]
  wire [15:0] n96_I_0_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_0_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_0_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_1_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_1_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_1_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_2_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_2_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_2_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_3_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_3_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_3_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_4_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_4_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_4_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_5_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_5_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_5_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_6_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_6_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_6_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_7_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_7_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_7_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_8_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_8_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_8_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_9_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_9_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_9_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_10_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_10_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_10_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_11_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_11_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_11_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_12_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_12_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_12_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_13_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_13_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_13_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_14_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_14_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_14_2; // @[Top.scala 140:21]
  wire [15:0] n96_I_15_0; // @[Top.scala 140:21]
  wire [15:0] n96_I_15_1; // @[Top.scala 140:21]
  wire [15:0] n96_I_15_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_0_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_0_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_0_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_1_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_1_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_1_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_2_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_2_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_2_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_3_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_3_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_3_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_4_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_4_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_4_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_5_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_5_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_5_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_6_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_6_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_6_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_7_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_7_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_7_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_8_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_8_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_8_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_9_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_9_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_9_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_10_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_10_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_10_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_11_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_11_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_11_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_12_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_12_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_12_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_13_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_13_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_13_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_14_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_14_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_14_2; // @[Top.scala 140:21]
  wire [15:0] n96_O_15_0; // @[Top.scala 140:21]
  wire [15:0] n96_O_15_1; // @[Top.scala 140:21]
  wire [15:0] n96_O_15_2; // @[Top.scala 140:21]
  wire  n97_valid_up; // @[Top.scala 143:21]
  wire  n97_valid_down; // @[Top.scala 143:21]
  wire [15:0] n97_I0_0_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_0_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_0_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_0_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_0_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_0_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_1_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_1_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_1_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_1_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_1_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_1_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_2_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_2_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_2_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_2_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_2_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_2_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_3_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_3_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_3_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_3_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_3_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_3_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_4_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_4_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_4_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_4_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_4_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_4_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_5_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_5_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_5_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_5_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_5_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_5_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_6_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_6_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_6_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_6_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_6_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_6_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_7_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_7_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_7_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_7_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_7_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_7_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_8_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_8_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_8_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_8_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_8_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_8_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_9_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_9_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_9_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_9_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_9_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_9_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_10_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_10_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_10_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_10_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_10_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_10_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_11_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_11_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_11_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_11_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_11_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_11_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_12_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_12_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_12_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_12_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_12_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_12_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_13_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_13_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_13_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_13_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_13_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_13_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_14_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_14_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_14_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_14_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_14_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_14_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_15_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_15_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_15_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I0_15_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I0_15_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I0_15_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_3_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_3_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_3_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_4_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_4_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_4_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_5_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_5_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_5_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_6_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_6_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_6_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_7_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_7_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_7_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_8_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_8_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_8_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_9_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_9_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_9_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_10_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_10_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_10_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_11_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_11_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_11_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_12_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_12_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_12_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_13_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_13_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_13_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_14_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_14_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_14_2; // @[Top.scala 143:21]
  wire [15:0] n97_I1_15_0; // @[Top.scala 143:21]
  wire [15:0] n97_I1_15_1; // @[Top.scala 143:21]
  wire [15:0] n97_I1_15_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_0_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_1_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_2_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_3_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_4_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_5_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_6_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_7_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_8_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_9_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_10_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_11_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_12_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_13_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_14_2_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_0_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_0_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_0_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_1_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_1_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_1_2; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_2_0; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_2_1; // @[Top.scala 143:21]
  wire [15:0] n97_O_15_2_2; // @[Top.scala 143:21]
  wire  n106_valid_up; // @[Top.scala 147:22]
  wire  n106_valid_down; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_1_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_2_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_3_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_4_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_5_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_6_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_7_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_8_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_9_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_10_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_11_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_12_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_13_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_14_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_I_15_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_0_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_1_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_2_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_3_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_4_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_5_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_6_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_7_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_8_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_9_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_10_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_11_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_12_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_13_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_14_0_2_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_0_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_0_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_0_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_1_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_1_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_1_2; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_2_0; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_2_1; // @[Top.scala 147:22]
  wire [15:0] n106_O_15_0_2_2; // @[Top.scala 147:22]
  wire  n113_valid_up; // @[Top.scala 150:22]
  wire  n113_valid_down; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_0_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_1_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_2_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_3_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_4_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_5_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_6_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_7_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_8_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_9_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_10_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_11_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_12_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_13_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_14_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_I_15_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_0_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_1_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_2_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_3_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_4_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_5_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_6_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_7_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_8_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_9_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_10_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_11_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_12_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_13_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_14_2_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_0_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_0_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_0_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_1_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_1_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_1_2; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_2_0; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_2_1; // @[Top.scala 150:22]
  wire [15:0] n113_O_15_2_2; // @[Top.scala 150:22]
  wire  n155_clock; // @[Top.scala 153:22]
  wire  n155_reset; // @[Top.scala 153:22]
  wire  n155_valid_up; // @[Top.scala 153:22]
  wire  n155_valid_down; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_0_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_1_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_2_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_3_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_4_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_5_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_6_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_7_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_8_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_9_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_10_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_11_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_12_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_13_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_14_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_0_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_0_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_1_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_1_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_1_2; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_2_0; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_2_1; // @[Top.scala 153:22]
  wire [15:0] n155_I_15_2_2; // @[Top.scala 153:22]
  wire [15:0] n155_O_0_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_1_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_2_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_3_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_4_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_5_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_6_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_7_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_8_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_9_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_10_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_11_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_12_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_13_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_14_0_0; // @[Top.scala 153:22]
  wire [15:0] n155_O_15_0_0; // @[Top.scala 153:22]
  wire  n156_valid_up; // @[Top.scala 156:22]
  wire  n156_valid_down; // @[Top.scala 156:22]
  wire [15:0] n156_I_0_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_1_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_2_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_3_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_4_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_5_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_6_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_7_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_8_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_9_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_10_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_11_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_12_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_13_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_14_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_I_15_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_0_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_1_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_2_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_3_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_4_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_5_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_6_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_7_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_8_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_9_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_10_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_11_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_12_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_13_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_14_0; // @[Top.scala 156:22]
  wire [15:0] n156_O_15_0; // @[Top.scala 156:22]
  wire  n157_valid_up; // @[Top.scala 159:22]
  wire  n157_valid_down; // @[Top.scala 159:22]
  wire [15:0] n157_I_0_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_1_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_2_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_3_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_4_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_5_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_6_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_7_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_8_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_9_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_10_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_11_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_12_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_13_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_14_0; // @[Top.scala 159:22]
  wire [15:0] n157_I_15_0; // @[Top.scala 159:22]
  wire [15:0] n157_O_0; // @[Top.scala 159:22]
  wire [15:0] n157_O_1; // @[Top.scala 159:22]
  wire [15:0] n157_O_2; // @[Top.scala 159:22]
  wire [15:0] n157_O_3; // @[Top.scala 159:22]
  wire [15:0] n157_O_4; // @[Top.scala 159:22]
  wire [15:0] n157_O_5; // @[Top.scala 159:22]
  wire [15:0] n157_O_6; // @[Top.scala 159:22]
  wire [15:0] n157_O_7; // @[Top.scala 159:22]
  wire [15:0] n157_O_8; // @[Top.scala 159:22]
  wire [15:0] n157_O_9; // @[Top.scala 159:22]
  wire [15:0] n157_O_10; // @[Top.scala 159:22]
  wire [15:0] n157_O_11; // @[Top.scala 159:22]
  wire [15:0] n157_O_12; // @[Top.scala 159:22]
  wire [15:0] n157_O_13; // @[Top.scala 159:22]
  wire [15:0] n157_O_14; // @[Top.scala 159:22]
  wire [15:0] n157_O_15; // @[Top.scala 159:22]
  wire  n158_clock; // @[Top.scala 162:22]
  wire  n158_reset; // @[Top.scala 162:22]
  wire  n158_valid_up; // @[Top.scala 162:22]
  wire  n158_valid_down; // @[Top.scala 162:22]
  wire [15:0] n158_I_0; // @[Top.scala 162:22]
  wire [15:0] n158_I_1; // @[Top.scala 162:22]
  wire [15:0] n158_I_2; // @[Top.scala 162:22]
  wire [15:0] n158_I_3; // @[Top.scala 162:22]
  wire [15:0] n158_I_4; // @[Top.scala 162:22]
  wire [15:0] n158_I_5; // @[Top.scala 162:22]
  wire [15:0] n158_I_6; // @[Top.scala 162:22]
  wire [15:0] n158_I_7; // @[Top.scala 162:22]
  wire [15:0] n158_I_8; // @[Top.scala 162:22]
  wire [15:0] n158_I_9; // @[Top.scala 162:22]
  wire [15:0] n158_I_10; // @[Top.scala 162:22]
  wire [15:0] n158_I_11; // @[Top.scala 162:22]
  wire [15:0] n158_I_12; // @[Top.scala 162:22]
  wire [15:0] n158_I_13; // @[Top.scala 162:22]
  wire [15:0] n158_I_14; // @[Top.scala 162:22]
  wire [15:0] n158_I_15; // @[Top.scala 162:22]
  wire [15:0] n158_O_0; // @[Top.scala 162:22]
  wire [15:0] n158_O_1; // @[Top.scala 162:22]
  wire [15:0] n158_O_2; // @[Top.scala 162:22]
  wire [15:0] n158_O_3; // @[Top.scala 162:22]
  wire [15:0] n158_O_4; // @[Top.scala 162:22]
  wire [15:0] n158_O_5; // @[Top.scala 162:22]
  wire [15:0] n158_O_6; // @[Top.scala 162:22]
  wire [15:0] n158_O_7; // @[Top.scala 162:22]
  wire [15:0] n158_O_8; // @[Top.scala 162:22]
  wire [15:0] n158_O_9; // @[Top.scala 162:22]
  wire [15:0] n158_O_10; // @[Top.scala 162:22]
  wire [15:0] n158_O_11; // @[Top.scala 162:22]
  wire [15:0] n158_O_12; // @[Top.scala 162:22]
  wire [15:0] n158_O_13; // @[Top.scala 162:22]
  wire [15:0] n158_O_14; // @[Top.scala 162:22]
  wire [15:0] n158_O_15; // @[Top.scala 162:22]
  wire  n159_clock; // @[Top.scala 165:22]
  wire  n159_reset; // @[Top.scala 165:22]
  wire  n159_valid_up; // @[Top.scala 165:22]
  wire  n159_valid_down; // @[Top.scala 165:22]
  wire [15:0] n159_I_0; // @[Top.scala 165:22]
  wire [15:0] n159_I_1; // @[Top.scala 165:22]
  wire [15:0] n159_I_2; // @[Top.scala 165:22]
  wire [15:0] n159_I_3; // @[Top.scala 165:22]
  wire [15:0] n159_I_4; // @[Top.scala 165:22]
  wire [15:0] n159_I_5; // @[Top.scala 165:22]
  wire [15:0] n159_I_6; // @[Top.scala 165:22]
  wire [15:0] n159_I_7; // @[Top.scala 165:22]
  wire [15:0] n159_I_8; // @[Top.scala 165:22]
  wire [15:0] n159_I_9; // @[Top.scala 165:22]
  wire [15:0] n159_I_10; // @[Top.scala 165:22]
  wire [15:0] n159_I_11; // @[Top.scala 165:22]
  wire [15:0] n159_I_12; // @[Top.scala 165:22]
  wire [15:0] n159_I_13; // @[Top.scala 165:22]
  wire [15:0] n159_I_14; // @[Top.scala 165:22]
  wire [15:0] n159_I_15; // @[Top.scala 165:22]
  wire [15:0] n159_O_0; // @[Top.scala 165:22]
  wire [15:0] n159_O_1; // @[Top.scala 165:22]
  wire [15:0] n159_O_2; // @[Top.scala 165:22]
  wire [15:0] n159_O_3; // @[Top.scala 165:22]
  wire [15:0] n159_O_4; // @[Top.scala 165:22]
  wire [15:0] n159_O_5; // @[Top.scala 165:22]
  wire [15:0] n159_O_6; // @[Top.scala 165:22]
  wire [15:0] n159_O_7; // @[Top.scala 165:22]
  wire [15:0] n159_O_8; // @[Top.scala 165:22]
  wire [15:0] n159_O_9; // @[Top.scala 165:22]
  wire [15:0] n159_O_10; // @[Top.scala 165:22]
  wire [15:0] n159_O_11; // @[Top.scala 165:22]
  wire [15:0] n159_O_12; // @[Top.scala 165:22]
  wire [15:0] n159_O_13; // @[Top.scala 165:22]
  wire [15:0] n159_O_14; // @[Top.scala 165:22]
  wire [15:0] n159_O_15; // @[Top.scala 165:22]
  wire  n160_clock; // @[Top.scala 168:22]
  wire  n160_reset; // @[Top.scala 168:22]
  wire  n160_valid_up; // @[Top.scala 168:22]
  wire  n160_valid_down; // @[Top.scala 168:22]
  wire [15:0] n160_I_0; // @[Top.scala 168:22]
  wire [15:0] n160_I_1; // @[Top.scala 168:22]
  wire [15:0] n160_I_2; // @[Top.scala 168:22]
  wire [15:0] n160_I_3; // @[Top.scala 168:22]
  wire [15:0] n160_I_4; // @[Top.scala 168:22]
  wire [15:0] n160_I_5; // @[Top.scala 168:22]
  wire [15:0] n160_I_6; // @[Top.scala 168:22]
  wire [15:0] n160_I_7; // @[Top.scala 168:22]
  wire [15:0] n160_I_8; // @[Top.scala 168:22]
  wire [15:0] n160_I_9; // @[Top.scala 168:22]
  wire [15:0] n160_I_10; // @[Top.scala 168:22]
  wire [15:0] n160_I_11; // @[Top.scala 168:22]
  wire [15:0] n160_I_12; // @[Top.scala 168:22]
  wire [15:0] n160_I_13; // @[Top.scala 168:22]
  wire [15:0] n160_I_14; // @[Top.scala 168:22]
  wire [15:0] n160_I_15; // @[Top.scala 168:22]
  wire [15:0] n160_O_0; // @[Top.scala 168:22]
  wire [15:0] n160_O_1; // @[Top.scala 168:22]
  wire [15:0] n160_O_2; // @[Top.scala 168:22]
  wire [15:0] n160_O_3; // @[Top.scala 168:22]
  wire [15:0] n160_O_4; // @[Top.scala 168:22]
  wire [15:0] n160_O_5; // @[Top.scala 168:22]
  wire [15:0] n160_O_6; // @[Top.scala 168:22]
  wire [15:0] n160_O_7; // @[Top.scala 168:22]
  wire [15:0] n160_O_8; // @[Top.scala 168:22]
  wire [15:0] n160_O_9; // @[Top.scala 168:22]
  wire [15:0] n160_O_10; // @[Top.scala 168:22]
  wire [15:0] n160_O_11; // @[Top.scala 168:22]
  wire [15:0] n160_O_12; // @[Top.scala 168:22]
  wire [15:0] n160_O_13; // @[Top.scala 168:22]
  wire [15:0] n160_O_14; // @[Top.scala 168:22]
  wire [15:0] n160_O_15; // @[Top.scala 168:22]
  FIFO n1 ( // @[Top.scala 46:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .I_8(n1_I_8),
    .I_9(n1_I_9),
    .I_10(n1_I_10),
    .I_11(n1_I_11),
    .I_12(n1_I_12),
    .I_13(n1_I_13),
    .I_14(n1_I_14),
    .I_15(n1_I_15),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7),
    .O_8(n1_O_8),
    .O_9(n1_O_9),
    .O_10(n1_O_10),
    .O_11(n1_O_11),
    .O_12(n1_O_12),
    .O_13(n1_O_13),
    .O_14(n1_O_14),
    .O_15(n1_O_15)
  );
  ShiftTS n2 ( // @[Top.scala 49:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .I_2(n2_I_2),
    .I_3(n2_I_3),
    .I_4(n2_I_4),
    .I_5(n2_I_5),
    .I_6(n2_I_6),
    .I_7(n2_I_7),
    .I_8(n2_I_8),
    .I_9(n2_I_9),
    .I_10(n2_I_10),
    .I_11(n2_I_11),
    .I_12(n2_I_12),
    .I_13(n2_I_13),
    .I_14(n2_I_14),
    .I_15(n2_I_15),
    .O_0(n2_O_0),
    .O_1(n2_O_1),
    .O_2(n2_O_2),
    .O_3(n2_O_3),
    .O_4(n2_O_4),
    .O_5(n2_O_5),
    .O_6(n2_O_6),
    .O_7(n2_O_7),
    .O_8(n2_O_8),
    .O_9(n2_O_9),
    .O_10(n2_O_10),
    .O_11(n2_O_11),
    .O_12(n2_O_12),
    .O_13(n2_O_13),
    .O_14(n2_O_14),
    .O_15(n2_O_15)
  );
  ShiftTS n3 ( // @[Top.scala 52:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .I_2(n3_I_2),
    .I_3(n3_I_3),
    .I_4(n3_I_4),
    .I_5(n3_I_5),
    .I_6(n3_I_6),
    .I_7(n3_I_7),
    .I_8(n3_I_8),
    .I_9(n3_I_9),
    .I_10(n3_I_10),
    .I_11(n3_I_11),
    .I_12(n3_I_12),
    .I_13(n3_I_13),
    .I_14(n3_I_14),
    .I_15(n3_I_15),
    .O_0(n3_O_0),
    .O_1(n3_O_1),
    .O_2(n3_O_2),
    .O_3(n3_O_3),
    .O_4(n3_O_4),
    .O_5(n3_O_5),
    .O_6(n3_O_6),
    .O_7(n3_O_7),
    .O_8(n3_O_8),
    .O_9(n3_O_9),
    .O_10(n3_O_10),
    .O_11(n3_O_11),
    .O_12(n3_O_12),
    .O_13(n3_O_13),
    .O_14(n3_O_14),
    .O_15(n3_O_15)
  );
  ShiftTS_2 n4 ( // @[Top.scala 55:20]
    .clock(n4_clock),
    .reset(n4_reset),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .I_2(n4_I_2),
    .I_3(n4_I_3),
    .I_4(n4_I_4),
    .I_5(n4_I_5),
    .I_6(n4_I_6),
    .I_7(n4_I_7),
    .I_8(n4_I_8),
    .I_9(n4_I_9),
    .I_10(n4_I_10),
    .I_11(n4_I_11),
    .I_12(n4_I_12),
    .I_13(n4_I_13),
    .I_14(n4_I_14),
    .I_15(n4_I_15),
    .O_0(n4_O_0),
    .O_1(n4_O_1),
    .O_2(n4_O_2),
    .O_3(n4_O_3),
    .O_4(n4_O_4),
    .O_5(n4_O_5),
    .O_6(n4_O_6),
    .O_7(n4_O_7),
    .O_8(n4_O_8),
    .O_9(n4_O_9),
    .O_10(n4_O_10),
    .O_11(n4_O_11),
    .O_12(n4_O_12),
    .O_13(n4_O_13),
    .O_14(n4_O_14),
    .O_15(n4_O_15)
  );
  ShiftTS_2 n5 ( // @[Top.scala 58:20]
    .clock(n5_clock),
    .reset(n5_reset),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .I_2(n5_I_2),
    .I_3(n5_I_3),
    .I_4(n5_I_4),
    .I_5(n5_I_5),
    .I_6(n5_I_6),
    .I_7(n5_I_7),
    .I_8(n5_I_8),
    .I_9(n5_I_9),
    .I_10(n5_I_10),
    .I_11(n5_I_11),
    .I_12(n5_I_12),
    .I_13(n5_I_13),
    .I_14(n5_I_14),
    .I_15(n5_I_15),
    .O_0(n5_O_0),
    .O_1(n5_O_1),
    .O_2(n5_O_2),
    .O_3(n5_O_3),
    .O_4(n5_O_4),
    .O_5(n5_O_5),
    .O_6(n5_O_6),
    .O_7(n5_O_7),
    .O_8(n5_O_8),
    .O_9(n5_O_9),
    .O_10(n5_O_10),
    .O_11(n5_O_11),
    .O_12(n5_O_12),
    .O_13(n5_O_13),
    .O_14(n5_O_14),
    .O_15(n5_O_15)
  );
  FIFO n6 ( // @[Top.scala 61:20]
    .clock(n6_clock),
    .reset(n6_reset),
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I_0(n6_I_0),
    .I_1(n6_I_1),
    .I_2(n6_I_2),
    .I_3(n6_I_3),
    .I_4(n6_I_4),
    .I_5(n6_I_5),
    .I_6(n6_I_6),
    .I_7(n6_I_7),
    .I_8(n6_I_8),
    .I_9(n6_I_9),
    .I_10(n6_I_10),
    .I_11(n6_I_11),
    .I_12(n6_I_12),
    .I_13(n6_I_13),
    .I_14(n6_I_14),
    .I_15(n6_I_15),
    .O_0(n6_O_0),
    .O_1(n6_O_1),
    .O_2(n6_O_2),
    .O_3(n6_O_3),
    .O_4(n6_O_4),
    .O_5(n6_O_5),
    .O_6(n6_O_6),
    .O_7(n6_O_7),
    .O_8(n6_O_8),
    .O_9(n6_O_9),
    .O_10(n6_O_10),
    .O_11(n6_O_11),
    .O_12(n6_O_12),
    .O_13(n6_O_13),
    .O_14(n6_O_14),
    .O_15(n6_O_15)
  );
  Map2T n7 ( // @[Top.scala 64:20]
    .valid_up(n7_valid_up),
    .valid_down(n7_valid_down),
    .I0_0(n7_I0_0),
    .I0_1(n7_I0_1),
    .I0_2(n7_I0_2),
    .I0_3(n7_I0_3),
    .I0_4(n7_I0_4),
    .I0_5(n7_I0_5),
    .I0_6(n7_I0_6),
    .I0_7(n7_I0_7),
    .I0_8(n7_I0_8),
    .I0_9(n7_I0_9),
    .I0_10(n7_I0_10),
    .I0_11(n7_I0_11),
    .I0_12(n7_I0_12),
    .I0_13(n7_I0_13),
    .I0_14(n7_I0_14),
    .I0_15(n7_I0_15),
    .I1_0(n7_I1_0),
    .I1_1(n7_I1_1),
    .I1_2(n7_I1_2),
    .I1_3(n7_I1_3),
    .I1_4(n7_I1_4),
    .I1_5(n7_I1_5),
    .I1_6(n7_I1_6),
    .I1_7(n7_I1_7),
    .I1_8(n7_I1_8),
    .I1_9(n7_I1_9),
    .I1_10(n7_I1_10),
    .I1_11(n7_I1_11),
    .I1_12(n7_I1_12),
    .I1_13(n7_I1_13),
    .I1_14(n7_I1_14),
    .I1_15(n7_I1_15),
    .O_0_0(n7_O_0_0),
    .O_0_1(n7_O_0_1),
    .O_1_0(n7_O_1_0),
    .O_1_1(n7_O_1_1),
    .O_2_0(n7_O_2_0),
    .O_2_1(n7_O_2_1),
    .O_3_0(n7_O_3_0),
    .O_3_1(n7_O_3_1),
    .O_4_0(n7_O_4_0),
    .O_4_1(n7_O_4_1),
    .O_5_0(n7_O_5_0),
    .O_5_1(n7_O_5_1),
    .O_6_0(n7_O_6_0),
    .O_6_1(n7_O_6_1),
    .O_7_0(n7_O_7_0),
    .O_7_1(n7_O_7_1),
    .O_8_0(n7_O_8_0),
    .O_8_1(n7_O_8_1),
    .O_9_0(n7_O_9_0),
    .O_9_1(n7_O_9_1),
    .O_10_0(n7_O_10_0),
    .O_10_1(n7_O_10_1),
    .O_11_0(n7_O_11_0),
    .O_11_1(n7_O_11_1),
    .O_12_0(n7_O_12_0),
    .O_12_1(n7_O_12_1),
    .O_13_0(n7_O_13_0),
    .O_13_1(n7_O_13_1),
    .O_14_0(n7_O_14_0),
    .O_14_1(n7_O_14_1),
    .O_15_0(n7_O_15_0),
    .O_15_1(n7_O_15_1)
  );
  FIFO_2 n14 ( // @[Top.scala 68:21]
    .clock(n14_clock),
    .reset(n14_reset),
    .valid_up(n14_valid_up),
    .valid_down(n14_valid_down),
    .I_0(n14_I_0),
    .I_1(n14_I_1),
    .I_2(n14_I_2),
    .I_3(n14_I_3),
    .I_4(n14_I_4),
    .I_5(n14_I_5),
    .I_6(n14_I_6),
    .I_7(n14_I_7),
    .I_8(n14_I_8),
    .I_9(n14_I_9),
    .I_10(n14_I_10),
    .I_11(n14_I_11),
    .I_12(n14_I_12),
    .I_13(n14_I_13),
    .I_14(n14_I_14),
    .I_15(n14_I_15),
    .O_0(n14_O_0),
    .O_1(n14_O_1),
    .O_2(n14_O_2),
    .O_3(n14_O_3),
    .O_4(n14_O_4),
    .O_5(n14_O_5),
    .O_6(n14_O_6),
    .O_7(n14_O_7),
    .O_8(n14_O_8),
    .O_9(n14_O_9),
    .O_10(n14_O_10),
    .O_11(n14_O_11),
    .O_12(n14_O_12),
    .O_13(n14_O_13),
    .O_14(n14_O_14),
    .O_15(n14_O_15)
  );
  Map2T_1 n15 ( // @[Top.scala 71:21]
    .valid_up(n15_valid_up),
    .valid_down(n15_valid_down),
    .I0_0_0(n15_I0_0_0),
    .I0_0_1(n15_I0_0_1),
    .I0_1_0(n15_I0_1_0),
    .I0_1_1(n15_I0_1_1),
    .I0_2_0(n15_I0_2_0),
    .I0_2_1(n15_I0_2_1),
    .I0_3_0(n15_I0_3_0),
    .I0_3_1(n15_I0_3_1),
    .I0_4_0(n15_I0_4_0),
    .I0_4_1(n15_I0_4_1),
    .I0_5_0(n15_I0_5_0),
    .I0_5_1(n15_I0_5_1),
    .I0_6_0(n15_I0_6_0),
    .I0_6_1(n15_I0_6_1),
    .I0_7_0(n15_I0_7_0),
    .I0_7_1(n15_I0_7_1),
    .I0_8_0(n15_I0_8_0),
    .I0_8_1(n15_I0_8_1),
    .I0_9_0(n15_I0_9_0),
    .I0_9_1(n15_I0_9_1),
    .I0_10_0(n15_I0_10_0),
    .I0_10_1(n15_I0_10_1),
    .I0_11_0(n15_I0_11_0),
    .I0_11_1(n15_I0_11_1),
    .I0_12_0(n15_I0_12_0),
    .I0_12_1(n15_I0_12_1),
    .I0_13_0(n15_I0_13_0),
    .I0_13_1(n15_I0_13_1),
    .I0_14_0(n15_I0_14_0),
    .I0_14_1(n15_I0_14_1),
    .I0_15_0(n15_I0_15_0),
    .I0_15_1(n15_I0_15_1),
    .I1_0(n15_I1_0),
    .I1_1(n15_I1_1),
    .I1_2(n15_I1_2),
    .I1_3(n15_I1_3),
    .I1_4(n15_I1_4),
    .I1_5(n15_I1_5),
    .I1_6(n15_I1_6),
    .I1_7(n15_I1_7),
    .I1_8(n15_I1_8),
    .I1_9(n15_I1_9),
    .I1_10(n15_I1_10),
    .I1_11(n15_I1_11),
    .I1_12(n15_I1_12),
    .I1_13(n15_I1_13),
    .I1_14(n15_I1_14),
    .I1_15(n15_I1_15),
    .O_0_0(n15_O_0_0),
    .O_0_1(n15_O_0_1),
    .O_0_2(n15_O_0_2),
    .O_1_0(n15_O_1_0),
    .O_1_1(n15_O_1_1),
    .O_1_2(n15_O_1_2),
    .O_2_0(n15_O_2_0),
    .O_2_1(n15_O_2_1),
    .O_2_2(n15_O_2_2),
    .O_3_0(n15_O_3_0),
    .O_3_1(n15_O_3_1),
    .O_3_2(n15_O_3_2),
    .O_4_0(n15_O_4_0),
    .O_4_1(n15_O_4_1),
    .O_4_2(n15_O_4_2),
    .O_5_0(n15_O_5_0),
    .O_5_1(n15_O_5_1),
    .O_5_2(n15_O_5_2),
    .O_6_0(n15_O_6_0),
    .O_6_1(n15_O_6_1),
    .O_6_2(n15_O_6_2),
    .O_7_0(n15_O_7_0),
    .O_7_1(n15_O_7_1),
    .O_7_2(n15_O_7_2),
    .O_8_0(n15_O_8_0),
    .O_8_1(n15_O_8_1),
    .O_8_2(n15_O_8_2),
    .O_9_0(n15_O_9_0),
    .O_9_1(n15_O_9_1),
    .O_9_2(n15_O_9_2),
    .O_10_0(n15_O_10_0),
    .O_10_1(n15_O_10_1),
    .O_10_2(n15_O_10_2),
    .O_11_0(n15_O_11_0),
    .O_11_1(n15_O_11_1),
    .O_11_2(n15_O_11_2),
    .O_12_0(n15_O_12_0),
    .O_12_1(n15_O_12_1),
    .O_12_2(n15_O_12_2),
    .O_13_0(n15_O_13_0),
    .O_13_1(n15_O_13_1),
    .O_13_2(n15_O_13_2),
    .O_14_0(n15_O_14_0),
    .O_14_1(n15_O_14_1),
    .O_14_2(n15_O_14_2),
    .O_15_0(n15_O_15_0),
    .O_15_1(n15_O_15_1),
    .O_15_2(n15_O_15_2)
  );
  MapT n24 ( // @[Top.scala 75:21]
    .valid_up(n24_valid_up),
    .valid_down(n24_valid_down),
    .I_0_0(n24_I_0_0),
    .I_0_1(n24_I_0_1),
    .I_0_2(n24_I_0_2),
    .I_1_0(n24_I_1_0),
    .I_1_1(n24_I_1_1),
    .I_1_2(n24_I_1_2),
    .I_2_0(n24_I_2_0),
    .I_2_1(n24_I_2_1),
    .I_2_2(n24_I_2_2),
    .I_3_0(n24_I_3_0),
    .I_3_1(n24_I_3_1),
    .I_3_2(n24_I_3_2),
    .I_4_0(n24_I_4_0),
    .I_4_1(n24_I_4_1),
    .I_4_2(n24_I_4_2),
    .I_5_0(n24_I_5_0),
    .I_5_1(n24_I_5_1),
    .I_5_2(n24_I_5_2),
    .I_6_0(n24_I_6_0),
    .I_6_1(n24_I_6_1),
    .I_6_2(n24_I_6_2),
    .I_7_0(n24_I_7_0),
    .I_7_1(n24_I_7_1),
    .I_7_2(n24_I_7_2),
    .I_8_0(n24_I_8_0),
    .I_8_1(n24_I_8_1),
    .I_8_2(n24_I_8_2),
    .I_9_0(n24_I_9_0),
    .I_9_1(n24_I_9_1),
    .I_9_2(n24_I_9_2),
    .I_10_0(n24_I_10_0),
    .I_10_1(n24_I_10_1),
    .I_10_2(n24_I_10_2),
    .I_11_0(n24_I_11_0),
    .I_11_1(n24_I_11_1),
    .I_11_2(n24_I_11_2),
    .I_12_0(n24_I_12_0),
    .I_12_1(n24_I_12_1),
    .I_12_2(n24_I_12_2),
    .I_13_0(n24_I_13_0),
    .I_13_1(n24_I_13_1),
    .I_13_2(n24_I_13_2),
    .I_14_0(n24_I_14_0),
    .I_14_1(n24_I_14_1),
    .I_14_2(n24_I_14_2),
    .I_15_0(n24_I_15_0),
    .I_15_1(n24_I_15_1),
    .I_15_2(n24_I_15_2),
    .O_0_0_0(n24_O_0_0_0),
    .O_0_0_1(n24_O_0_0_1),
    .O_0_0_2(n24_O_0_0_2),
    .O_1_0_0(n24_O_1_0_0),
    .O_1_0_1(n24_O_1_0_1),
    .O_1_0_2(n24_O_1_0_2),
    .O_2_0_0(n24_O_2_0_0),
    .O_2_0_1(n24_O_2_0_1),
    .O_2_0_2(n24_O_2_0_2),
    .O_3_0_0(n24_O_3_0_0),
    .O_3_0_1(n24_O_3_0_1),
    .O_3_0_2(n24_O_3_0_2),
    .O_4_0_0(n24_O_4_0_0),
    .O_4_0_1(n24_O_4_0_1),
    .O_4_0_2(n24_O_4_0_2),
    .O_5_0_0(n24_O_5_0_0),
    .O_5_0_1(n24_O_5_0_1),
    .O_5_0_2(n24_O_5_0_2),
    .O_6_0_0(n24_O_6_0_0),
    .O_6_0_1(n24_O_6_0_1),
    .O_6_0_2(n24_O_6_0_2),
    .O_7_0_0(n24_O_7_0_0),
    .O_7_0_1(n24_O_7_0_1),
    .O_7_0_2(n24_O_7_0_2),
    .O_8_0_0(n24_O_8_0_0),
    .O_8_0_1(n24_O_8_0_1),
    .O_8_0_2(n24_O_8_0_2),
    .O_9_0_0(n24_O_9_0_0),
    .O_9_0_1(n24_O_9_0_1),
    .O_9_0_2(n24_O_9_0_2),
    .O_10_0_0(n24_O_10_0_0),
    .O_10_0_1(n24_O_10_0_1),
    .O_10_0_2(n24_O_10_0_2),
    .O_11_0_0(n24_O_11_0_0),
    .O_11_0_1(n24_O_11_0_1),
    .O_11_0_2(n24_O_11_0_2),
    .O_12_0_0(n24_O_12_0_0),
    .O_12_0_1(n24_O_12_0_1),
    .O_12_0_2(n24_O_12_0_2),
    .O_13_0_0(n24_O_13_0_0),
    .O_13_0_1(n24_O_13_0_1),
    .O_13_0_2(n24_O_13_0_2),
    .O_14_0_0(n24_O_14_0_0),
    .O_14_0_1(n24_O_14_0_1),
    .O_14_0_2(n24_O_14_0_2),
    .O_15_0_0(n24_O_15_0_0),
    .O_15_0_1(n24_O_15_0_1),
    .O_15_0_2(n24_O_15_0_2)
  );
  MapT_1 n31 ( // @[Top.scala 78:21]
    .valid_up(n31_valid_up),
    .valid_down(n31_valid_down),
    .I_0_0_0(n31_I_0_0_0),
    .I_0_0_1(n31_I_0_0_1),
    .I_0_0_2(n31_I_0_0_2),
    .I_1_0_0(n31_I_1_0_0),
    .I_1_0_1(n31_I_1_0_1),
    .I_1_0_2(n31_I_1_0_2),
    .I_2_0_0(n31_I_2_0_0),
    .I_2_0_1(n31_I_2_0_1),
    .I_2_0_2(n31_I_2_0_2),
    .I_3_0_0(n31_I_3_0_0),
    .I_3_0_1(n31_I_3_0_1),
    .I_3_0_2(n31_I_3_0_2),
    .I_4_0_0(n31_I_4_0_0),
    .I_4_0_1(n31_I_4_0_1),
    .I_4_0_2(n31_I_4_0_2),
    .I_5_0_0(n31_I_5_0_0),
    .I_5_0_1(n31_I_5_0_1),
    .I_5_0_2(n31_I_5_0_2),
    .I_6_0_0(n31_I_6_0_0),
    .I_6_0_1(n31_I_6_0_1),
    .I_6_0_2(n31_I_6_0_2),
    .I_7_0_0(n31_I_7_0_0),
    .I_7_0_1(n31_I_7_0_1),
    .I_7_0_2(n31_I_7_0_2),
    .I_8_0_0(n31_I_8_0_0),
    .I_8_0_1(n31_I_8_0_1),
    .I_8_0_2(n31_I_8_0_2),
    .I_9_0_0(n31_I_9_0_0),
    .I_9_0_1(n31_I_9_0_1),
    .I_9_0_2(n31_I_9_0_2),
    .I_10_0_0(n31_I_10_0_0),
    .I_10_0_1(n31_I_10_0_1),
    .I_10_0_2(n31_I_10_0_2),
    .I_11_0_0(n31_I_11_0_0),
    .I_11_0_1(n31_I_11_0_1),
    .I_11_0_2(n31_I_11_0_2),
    .I_12_0_0(n31_I_12_0_0),
    .I_12_0_1(n31_I_12_0_1),
    .I_12_0_2(n31_I_12_0_2),
    .I_13_0_0(n31_I_13_0_0),
    .I_13_0_1(n31_I_13_0_1),
    .I_13_0_2(n31_I_13_0_2),
    .I_14_0_0(n31_I_14_0_0),
    .I_14_0_1(n31_I_14_0_1),
    .I_14_0_2(n31_I_14_0_2),
    .I_15_0_0(n31_I_15_0_0),
    .I_15_0_1(n31_I_15_0_1),
    .I_15_0_2(n31_I_15_0_2),
    .O_0_0(n31_O_0_0),
    .O_0_1(n31_O_0_1),
    .O_0_2(n31_O_0_2),
    .O_1_0(n31_O_1_0),
    .O_1_1(n31_O_1_1),
    .O_1_2(n31_O_1_2),
    .O_2_0(n31_O_2_0),
    .O_2_1(n31_O_2_1),
    .O_2_2(n31_O_2_2),
    .O_3_0(n31_O_3_0),
    .O_3_1(n31_O_3_1),
    .O_3_2(n31_O_3_2),
    .O_4_0(n31_O_4_0),
    .O_4_1(n31_O_4_1),
    .O_4_2(n31_O_4_2),
    .O_5_0(n31_O_5_0),
    .O_5_1(n31_O_5_1),
    .O_5_2(n31_O_5_2),
    .O_6_0(n31_O_6_0),
    .O_6_1(n31_O_6_1),
    .O_6_2(n31_O_6_2),
    .O_7_0(n31_O_7_0),
    .O_7_1(n31_O_7_1),
    .O_7_2(n31_O_7_2),
    .O_8_0(n31_O_8_0),
    .O_8_1(n31_O_8_1),
    .O_8_2(n31_O_8_2),
    .O_9_0(n31_O_9_0),
    .O_9_1(n31_O_9_1),
    .O_9_2(n31_O_9_2),
    .O_10_0(n31_O_10_0),
    .O_10_1(n31_O_10_1),
    .O_10_2(n31_O_10_2),
    .O_11_0(n31_O_11_0),
    .O_11_1(n31_O_11_1),
    .O_11_2(n31_O_11_2),
    .O_12_0(n31_O_12_0),
    .O_12_1(n31_O_12_1),
    .O_12_2(n31_O_12_2),
    .O_13_0(n31_O_13_0),
    .O_13_1(n31_O_13_1),
    .O_13_2(n31_O_13_2),
    .O_14_0(n31_O_14_0),
    .O_14_1(n31_O_14_1),
    .O_14_2(n31_O_14_2),
    .O_15_0(n31_O_15_0),
    .O_15_1(n31_O_15_1),
    .O_15_2(n31_O_15_2)
  );
  ShiftTS_2 n32 ( // @[Top.scala 81:21]
    .clock(n32_clock),
    .reset(n32_reset),
    .valid_up(n32_valid_up),
    .valid_down(n32_valid_down),
    .I_0(n32_I_0),
    .I_1(n32_I_1),
    .I_2(n32_I_2),
    .I_3(n32_I_3),
    .I_4(n32_I_4),
    .I_5(n32_I_5),
    .I_6(n32_I_6),
    .I_7(n32_I_7),
    .I_8(n32_I_8),
    .I_9(n32_I_9),
    .I_10(n32_I_10),
    .I_11(n32_I_11),
    .I_12(n32_I_12),
    .I_13(n32_I_13),
    .I_14(n32_I_14),
    .I_15(n32_I_15),
    .O_0(n32_O_0),
    .O_1(n32_O_1),
    .O_2(n32_O_2),
    .O_3(n32_O_3),
    .O_4(n32_O_4),
    .O_5(n32_O_5),
    .O_6(n32_O_6),
    .O_7(n32_O_7),
    .O_8(n32_O_8),
    .O_9(n32_O_9),
    .O_10(n32_O_10),
    .O_11(n32_O_11),
    .O_12(n32_O_12),
    .O_13(n32_O_13),
    .O_14(n32_O_14),
    .O_15(n32_O_15)
  );
  ShiftTS_2 n33 ( // @[Top.scala 84:21]
    .clock(n33_clock),
    .reset(n33_reset),
    .valid_up(n33_valid_up),
    .valid_down(n33_valid_down),
    .I_0(n33_I_0),
    .I_1(n33_I_1),
    .I_2(n33_I_2),
    .I_3(n33_I_3),
    .I_4(n33_I_4),
    .I_5(n33_I_5),
    .I_6(n33_I_6),
    .I_7(n33_I_7),
    .I_8(n33_I_8),
    .I_9(n33_I_9),
    .I_10(n33_I_10),
    .I_11(n33_I_11),
    .I_12(n33_I_12),
    .I_13(n33_I_13),
    .I_14(n33_I_14),
    .I_15(n33_I_15),
    .O_0(n33_O_0),
    .O_1(n33_O_1),
    .O_2(n33_O_2),
    .O_3(n33_O_3),
    .O_4(n33_O_4),
    .O_5(n33_O_5),
    .O_6(n33_O_6),
    .O_7(n33_O_7),
    .O_8(n33_O_8),
    .O_9(n33_O_9),
    .O_10(n33_O_10),
    .O_11(n33_O_11),
    .O_12(n33_O_12),
    .O_13(n33_O_13),
    .O_14(n33_O_14),
    .O_15(n33_O_15)
  );
  FIFO n34 ( // @[Top.scala 87:21]
    .clock(n34_clock),
    .reset(n34_reset),
    .valid_up(n34_valid_up),
    .valid_down(n34_valid_down),
    .I_0(n34_I_0),
    .I_1(n34_I_1),
    .I_2(n34_I_2),
    .I_3(n34_I_3),
    .I_4(n34_I_4),
    .I_5(n34_I_5),
    .I_6(n34_I_6),
    .I_7(n34_I_7),
    .I_8(n34_I_8),
    .I_9(n34_I_9),
    .I_10(n34_I_10),
    .I_11(n34_I_11),
    .I_12(n34_I_12),
    .I_13(n34_I_13),
    .I_14(n34_I_14),
    .I_15(n34_I_15),
    .O_0(n34_O_0),
    .O_1(n34_O_1),
    .O_2(n34_O_2),
    .O_3(n34_O_3),
    .O_4(n34_O_4),
    .O_5(n34_O_5),
    .O_6(n34_O_6),
    .O_7(n34_O_7),
    .O_8(n34_O_8),
    .O_9(n34_O_9),
    .O_10(n34_O_10),
    .O_11(n34_O_11),
    .O_12(n34_O_12),
    .O_13(n34_O_13),
    .O_14(n34_O_14),
    .O_15(n34_O_15)
  );
  Map2T n35 ( // @[Top.scala 90:21]
    .valid_up(n35_valid_up),
    .valid_down(n35_valid_down),
    .I0_0(n35_I0_0),
    .I0_1(n35_I0_1),
    .I0_2(n35_I0_2),
    .I0_3(n35_I0_3),
    .I0_4(n35_I0_4),
    .I0_5(n35_I0_5),
    .I0_6(n35_I0_6),
    .I0_7(n35_I0_7),
    .I0_8(n35_I0_8),
    .I0_9(n35_I0_9),
    .I0_10(n35_I0_10),
    .I0_11(n35_I0_11),
    .I0_12(n35_I0_12),
    .I0_13(n35_I0_13),
    .I0_14(n35_I0_14),
    .I0_15(n35_I0_15),
    .I1_0(n35_I1_0),
    .I1_1(n35_I1_1),
    .I1_2(n35_I1_2),
    .I1_3(n35_I1_3),
    .I1_4(n35_I1_4),
    .I1_5(n35_I1_5),
    .I1_6(n35_I1_6),
    .I1_7(n35_I1_7),
    .I1_8(n35_I1_8),
    .I1_9(n35_I1_9),
    .I1_10(n35_I1_10),
    .I1_11(n35_I1_11),
    .I1_12(n35_I1_12),
    .I1_13(n35_I1_13),
    .I1_14(n35_I1_14),
    .I1_15(n35_I1_15),
    .O_0_0(n35_O_0_0),
    .O_0_1(n35_O_0_1),
    .O_1_0(n35_O_1_0),
    .O_1_1(n35_O_1_1),
    .O_2_0(n35_O_2_0),
    .O_2_1(n35_O_2_1),
    .O_3_0(n35_O_3_0),
    .O_3_1(n35_O_3_1),
    .O_4_0(n35_O_4_0),
    .O_4_1(n35_O_4_1),
    .O_5_0(n35_O_5_0),
    .O_5_1(n35_O_5_1),
    .O_6_0(n35_O_6_0),
    .O_6_1(n35_O_6_1),
    .O_7_0(n35_O_7_0),
    .O_7_1(n35_O_7_1),
    .O_8_0(n35_O_8_0),
    .O_8_1(n35_O_8_1),
    .O_9_0(n35_O_9_0),
    .O_9_1(n35_O_9_1),
    .O_10_0(n35_O_10_0),
    .O_10_1(n35_O_10_1),
    .O_11_0(n35_O_11_0),
    .O_11_1(n35_O_11_1),
    .O_12_0(n35_O_12_0),
    .O_12_1(n35_O_12_1),
    .O_13_0(n35_O_13_0),
    .O_13_1(n35_O_13_1),
    .O_14_0(n35_O_14_0),
    .O_14_1(n35_O_14_1),
    .O_15_0(n35_O_15_0),
    .O_15_1(n35_O_15_1)
  );
  FIFO_2 n42 ( // @[Top.scala 94:21]
    .clock(n42_clock),
    .reset(n42_reset),
    .valid_up(n42_valid_up),
    .valid_down(n42_valid_down),
    .I_0(n42_I_0),
    .I_1(n42_I_1),
    .I_2(n42_I_2),
    .I_3(n42_I_3),
    .I_4(n42_I_4),
    .I_5(n42_I_5),
    .I_6(n42_I_6),
    .I_7(n42_I_7),
    .I_8(n42_I_8),
    .I_9(n42_I_9),
    .I_10(n42_I_10),
    .I_11(n42_I_11),
    .I_12(n42_I_12),
    .I_13(n42_I_13),
    .I_14(n42_I_14),
    .I_15(n42_I_15),
    .O_0(n42_O_0),
    .O_1(n42_O_1),
    .O_2(n42_O_2),
    .O_3(n42_O_3),
    .O_4(n42_O_4),
    .O_5(n42_O_5),
    .O_6(n42_O_6),
    .O_7(n42_O_7),
    .O_8(n42_O_8),
    .O_9(n42_O_9),
    .O_10(n42_O_10),
    .O_11(n42_O_11),
    .O_12(n42_O_12),
    .O_13(n42_O_13),
    .O_14(n42_O_14),
    .O_15(n42_O_15)
  );
  Map2T_1 n43 ( // @[Top.scala 97:21]
    .valid_up(n43_valid_up),
    .valid_down(n43_valid_down),
    .I0_0_0(n43_I0_0_0),
    .I0_0_1(n43_I0_0_1),
    .I0_1_0(n43_I0_1_0),
    .I0_1_1(n43_I0_1_1),
    .I0_2_0(n43_I0_2_0),
    .I0_2_1(n43_I0_2_1),
    .I0_3_0(n43_I0_3_0),
    .I0_3_1(n43_I0_3_1),
    .I0_4_0(n43_I0_4_0),
    .I0_4_1(n43_I0_4_1),
    .I0_5_0(n43_I0_5_0),
    .I0_5_1(n43_I0_5_1),
    .I0_6_0(n43_I0_6_0),
    .I0_6_1(n43_I0_6_1),
    .I0_7_0(n43_I0_7_0),
    .I0_7_1(n43_I0_7_1),
    .I0_8_0(n43_I0_8_0),
    .I0_8_1(n43_I0_8_1),
    .I0_9_0(n43_I0_9_0),
    .I0_9_1(n43_I0_9_1),
    .I0_10_0(n43_I0_10_0),
    .I0_10_1(n43_I0_10_1),
    .I0_11_0(n43_I0_11_0),
    .I0_11_1(n43_I0_11_1),
    .I0_12_0(n43_I0_12_0),
    .I0_12_1(n43_I0_12_1),
    .I0_13_0(n43_I0_13_0),
    .I0_13_1(n43_I0_13_1),
    .I0_14_0(n43_I0_14_0),
    .I0_14_1(n43_I0_14_1),
    .I0_15_0(n43_I0_15_0),
    .I0_15_1(n43_I0_15_1),
    .I1_0(n43_I1_0),
    .I1_1(n43_I1_1),
    .I1_2(n43_I1_2),
    .I1_3(n43_I1_3),
    .I1_4(n43_I1_4),
    .I1_5(n43_I1_5),
    .I1_6(n43_I1_6),
    .I1_7(n43_I1_7),
    .I1_8(n43_I1_8),
    .I1_9(n43_I1_9),
    .I1_10(n43_I1_10),
    .I1_11(n43_I1_11),
    .I1_12(n43_I1_12),
    .I1_13(n43_I1_13),
    .I1_14(n43_I1_14),
    .I1_15(n43_I1_15),
    .O_0_0(n43_O_0_0),
    .O_0_1(n43_O_0_1),
    .O_0_2(n43_O_0_2),
    .O_1_0(n43_O_1_0),
    .O_1_1(n43_O_1_1),
    .O_1_2(n43_O_1_2),
    .O_2_0(n43_O_2_0),
    .O_2_1(n43_O_2_1),
    .O_2_2(n43_O_2_2),
    .O_3_0(n43_O_3_0),
    .O_3_1(n43_O_3_1),
    .O_3_2(n43_O_3_2),
    .O_4_0(n43_O_4_0),
    .O_4_1(n43_O_4_1),
    .O_4_2(n43_O_4_2),
    .O_5_0(n43_O_5_0),
    .O_5_1(n43_O_5_1),
    .O_5_2(n43_O_5_2),
    .O_6_0(n43_O_6_0),
    .O_6_1(n43_O_6_1),
    .O_6_2(n43_O_6_2),
    .O_7_0(n43_O_7_0),
    .O_7_1(n43_O_7_1),
    .O_7_2(n43_O_7_2),
    .O_8_0(n43_O_8_0),
    .O_8_1(n43_O_8_1),
    .O_8_2(n43_O_8_2),
    .O_9_0(n43_O_9_0),
    .O_9_1(n43_O_9_1),
    .O_9_2(n43_O_9_2),
    .O_10_0(n43_O_10_0),
    .O_10_1(n43_O_10_1),
    .O_10_2(n43_O_10_2),
    .O_11_0(n43_O_11_0),
    .O_11_1(n43_O_11_1),
    .O_11_2(n43_O_11_2),
    .O_12_0(n43_O_12_0),
    .O_12_1(n43_O_12_1),
    .O_12_2(n43_O_12_2),
    .O_13_0(n43_O_13_0),
    .O_13_1(n43_O_13_1),
    .O_13_2(n43_O_13_2),
    .O_14_0(n43_O_14_0),
    .O_14_1(n43_O_14_1),
    .O_14_2(n43_O_14_2),
    .O_15_0(n43_O_15_0),
    .O_15_1(n43_O_15_1),
    .O_15_2(n43_O_15_2)
  );
  MapT n52 ( // @[Top.scala 101:21]
    .valid_up(n52_valid_up),
    .valid_down(n52_valid_down),
    .I_0_0(n52_I_0_0),
    .I_0_1(n52_I_0_1),
    .I_0_2(n52_I_0_2),
    .I_1_0(n52_I_1_0),
    .I_1_1(n52_I_1_1),
    .I_1_2(n52_I_1_2),
    .I_2_0(n52_I_2_0),
    .I_2_1(n52_I_2_1),
    .I_2_2(n52_I_2_2),
    .I_3_0(n52_I_3_0),
    .I_3_1(n52_I_3_1),
    .I_3_2(n52_I_3_2),
    .I_4_0(n52_I_4_0),
    .I_4_1(n52_I_4_1),
    .I_4_2(n52_I_4_2),
    .I_5_0(n52_I_5_0),
    .I_5_1(n52_I_5_1),
    .I_5_2(n52_I_5_2),
    .I_6_0(n52_I_6_0),
    .I_6_1(n52_I_6_1),
    .I_6_2(n52_I_6_2),
    .I_7_0(n52_I_7_0),
    .I_7_1(n52_I_7_1),
    .I_7_2(n52_I_7_2),
    .I_8_0(n52_I_8_0),
    .I_8_1(n52_I_8_1),
    .I_8_2(n52_I_8_2),
    .I_9_0(n52_I_9_0),
    .I_9_1(n52_I_9_1),
    .I_9_2(n52_I_9_2),
    .I_10_0(n52_I_10_0),
    .I_10_1(n52_I_10_1),
    .I_10_2(n52_I_10_2),
    .I_11_0(n52_I_11_0),
    .I_11_1(n52_I_11_1),
    .I_11_2(n52_I_11_2),
    .I_12_0(n52_I_12_0),
    .I_12_1(n52_I_12_1),
    .I_12_2(n52_I_12_2),
    .I_13_0(n52_I_13_0),
    .I_13_1(n52_I_13_1),
    .I_13_2(n52_I_13_2),
    .I_14_0(n52_I_14_0),
    .I_14_1(n52_I_14_1),
    .I_14_2(n52_I_14_2),
    .I_15_0(n52_I_15_0),
    .I_15_1(n52_I_15_1),
    .I_15_2(n52_I_15_2),
    .O_0_0_0(n52_O_0_0_0),
    .O_0_0_1(n52_O_0_0_1),
    .O_0_0_2(n52_O_0_0_2),
    .O_1_0_0(n52_O_1_0_0),
    .O_1_0_1(n52_O_1_0_1),
    .O_1_0_2(n52_O_1_0_2),
    .O_2_0_0(n52_O_2_0_0),
    .O_2_0_1(n52_O_2_0_1),
    .O_2_0_2(n52_O_2_0_2),
    .O_3_0_0(n52_O_3_0_0),
    .O_3_0_1(n52_O_3_0_1),
    .O_3_0_2(n52_O_3_0_2),
    .O_4_0_0(n52_O_4_0_0),
    .O_4_0_1(n52_O_4_0_1),
    .O_4_0_2(n52_O_4_0_2),
    .O_5_0_0(n52_O_5_0_0),
    .O_5_0_1(n52_O_5_0_1),
    .O_5_0_2(n52_O_5_0_2),
    .O_6_0_0(n52_O_6_0_0),
    .O_6_0_1(n52_O_6_0_1),
    .O_6_0_2(n52_O_6_0_2),
    .O_7_0_0(n52_O_7_0_0),
    .O_7_0_1(n52_O_7_0_1),
    .O_7_0_2(n52_O_7_0_2),
    .O_8_0_0(n52_O_8_0_0),
    .O_8_0_1(n52_O_8_0_1),
    .O_8_0_2(n52_O_8_0_2),
    .O_9_0_0(n52_O_9_0_0),
    .O_9_0_1(n52_O_9_0_1),
    .O_9_0_2(n52_O_9_0_2),
    .O_10_0_0(n52_O_10_0_0),
    .O_10_0_1(n52_O_10_0_1),
    .O_10_0_2(n52_O_10_0_2),
    .O_11_0_0(n52_O_11_0_0),
    .O_11_0_1(n52_O_11_0_1),
    .O_11_0_2(n52_O_11_0_2),
    .O_12_0_0(n52_O_12_0_0),
    .O_12_0_1(n52_O_12_0_1),
    .O_12_0_2(n52_O_12_0_2),
    .O_13_0_0(n52_O_13_0_0),
    .O_13_0_1(n52_O_13_0_1),
    .O_13_0_2(n52_O_13_0_2),
    .O_14_0_0(n52_O_14_0_0),
    .O_14_0_1(n52_O_14_0_1),
    .O_14_0_2(n52_O_14_0_2),
    .O_15_0_0(n52_O_15_0_0),
    .O_15_0_1(n52_O_15_0_1),
    .O_15_0_2(n52_O_15_0_2)
  );
  MapT_1 n59 ( // @[Top.scala 104:21]
    .valid_up(n59_valid_up),
    .valid_down(n59_valid_down),
    .I_0_0_0(n59_I_0_0_0),
    .I_0_0_1(n59_I_0_0_1),
    .I_0_0_2(n59_I_0_0_2),
    .I_1_0_0(n59_I_1_0_0),
    .I_1_0_1(n59_I_1_0_1),
    .I_1_0_2(n59_I_1_0_2),
    .I_2_0_0(n59_I_2_0_0),
    .I_2_0_1(n59_I_2_0_1),
    .I_2_0_2(n59_I_2_0_2),
    .I_3_0_0(n59_I_3_0_0),
    .I_3_0_1(n59_I_3_0_1),
    .I_3_0_2(n59_I_3_0_2),
    .I_4_0_0(n59_I_4_0_0),
    .I_4_0_1(n59_I_4_0_1),
    .I_4_0_2(n59_I_4_0_2),
    .I_5_0_0(n59_I_5_0_0),
    .I_5_0_1(n59_I_5_0_1),
    .I_5_0_2(n59_I_5_0_2),
    .I_6_0_0(n59_I_6_0_0),
    .I_6_0_1(n59_I_6_0_1),
    .I_6_0_2(n59_I_6_0_2),
    .I_7_0_0(n59_I_7_0_0),
    .I_7_0_1(n59_I_7_0_1),
    .I_7_0_2(n59_I_7_0_2),
    .I_8_0_0(n59_I_8_0_0),
    .I_8_0_1(n59_I_8_0_1),
    .I_8_0_2(n59_I_8_0_2),
    .I_9_0_0(n59_I_9_0_0),
    .I_9_0_1(n59_I_9_0_1),
    .I_9_0_2(n59_I_9_0_2),
    .I_10_0_0(n59_I_10_0_0),
    .I_10_0_1(n59_I_10_0_1),
    .I_10_0_2(n59_I_10_0_2),
    .I_11_0_0(n59_I_11_0_0),
    .I_11_0_1(n59_I_11_0_1),
    .I_11_0_2(n59_I_11_0_2),
    .I_12_0_0(n59_I_12_0_0),
    .I_12_0_1(n59_I_12_0_1),
    .I_12_0_2(n59_I_12_0_2),
    .I_13_0_0(n59_I_13_0_0),
    .I_13_0_1(n59_I_13_0_1),
    .I_13_0_2(n59_I_13_0_2),
    .I_14_0_0(n59_I_14_0_0),
    .I_14_0_1(n59_I_14_0_1),
    .I_14_0_2(n59_I_14_0_2),
    .I_15_0_0(n59_I_15_0_0),
    .I_15_0_1(n59_I_15_0_1),
    .I_15_0_2(n59_I_15_0_2),
    .O_0_0(n59_O_0_0),
    .O_0_1(n59_O_0_1),
    .O_0_2(n59_O_0_2),
    .O_1_0(n59_O_1_0),
    .O_1_1(n59_O_1_1),
    .O_1_2(n59_O_1_2),
    .O_2_0(n59_O_2_0),
    .O_2_1(n59_O_2_1),
    .O_2_2(n59_O_2_2),
    .O_3_0(n59_O_3_0),
    .O_3_1(n59_O_3_1),
    .O_3_2(n59_O_3_2),
    .O_4_0(n59_O_4_0),
    .O_4_1(n59_O_4_1),
    .O_4_2(n59_O_4_2),
    .O_5_0(n59_O_5_0),
    .O_5_1(n59_O_5_1),
    .O_5_2(n59_O_5_2),
    .O_6_0(n59_O_6_0),
    .O_6_1(n59_O_6_1),
    .O_6_2(n59_O_6_2),
    .O_7_0(n59_O_7_0),
    .O_7_1(n59_O_7_1),
    .O_7_2(n59_O_7_2),
    .O_8_0(n59_O_8_0),
    .O_8_1(n59_O_8_1),
    .O_8_2(n59_O_8_2),
    .O_9_0(n59_O_9_0),
    .O_9_1(n59_O_9_1),
    .O_9_2(n59_O_9_2),
    .O_10_0(n59_O_10_0),
    .O_10_1(n59_O_10_1),
    .O_10_2(n59_O_10_2),
    .O_11_0(n59_O_11_0),
    .O_11_1(n59_O_11_1),
    .O_11_2(n59_O_11_2),
    .O_12_0(n59_O_12_0),
    .O_12_1(n59_O_12_1),
    .O_12_2(n59_O_12_2),
    .O_13_0(n59_O_13_0),
    .O_13_1(n59_O_13_1),
    .O_13_2(n59_O_13_2),
    .O_14_0(n59_O_14_0),
    .O_14_1(n59_O_14_1),
    .O_14_2(n59_O_14_2),
    .O_15_0(n59_O_15_0),
    .O_15_1(n59_O_15_1),
    .O_15_2(n59_O_15_2)
  );
  FIFO_5 n60 ( // @[Top.scala 107:21]
    .clock(n60_clock),
    .reset(n60_reset),
    .valid_up(n60_valid_up),
    .valid_down(n60_valid_down),
    .I_0_0(n60_I_0_0),
    .I_0_1(n60_I_0_1),
    .I_0_2(n60_I_0_2),
    .I_1_0(n60_I_1_0),
    .I_1_1(n60_I_1_1),
    .I_1_2(n60_I_1_2),
    .I_2_0(n60_I_2_0),
    .I_2_1(n60_I_2_1),
    .I_2_2(n60_I_2_2),
    .I_3_0(n60_I_3_0),
    .I_3_1(n60_I_3_1),
    .I_3_2(n60_I_3_2),
    .I_4_0(n60_I_4_0),
    .I_4_1(n60_I_4_1),
    .I_4_2(n60_I_4_2),
    .I_5_0(n60_I_5_0),
    .I_5_1(n60_I_5_1),
    .I_5_2(n60_I_5_2),
    .I_6_0(n60_I_6_0),
    .I_6_1(n60_I_6_1),
    .I_6_2(n60_I_6_2),
    .I_7_0(n60_I_7_0),
    .I_7_1(n60_I_7_1),
    .I_7_2(n60_I_7_2),
    .I_8_0(n60_I_8_0),
    .I_8_1(n60_I_8_1),
    .I_8_2(n60_I_8_2),
    .I_9_0(n60_I_9_0),
    .I_9_1(n60_I_9_1),
    .I_9_2(n60_I_9_2),
    .I_10_0(n60_I_10_0),
    .I_10_1(n60_I_10_1),
    .I_10_2(n60_I_10_2),
    .I_11_0(n60_I_11_0),
    .I_11_1(n60_I_11_1),
    .I_11_2(n60_I_11_2),
    .I_12_0(n60_I_12_0),
    .I_12_1(n60_I_12_1),
    .I_12_2(n60_I_12_2),
    .I_13_0(n60_I_13_0),
    .I_13_1(n60_I_13_1),
    .I_13_2(n60_I_13_2),
    .I_14_0(n60_I_14_0),
    .I_14_1(n60_I_14_1),
    .I_14_2(n60_I_14_2),
    .I_15_0(n60_I_15_0),
    .I_15_1(n60_I_15_1),
    .I_15_2(n60_I_15_2),
    .O_0_0(n60_O_0_0),
    .O_0_1(n60_O_0_1),
    .O_0_2(n60_O_0_2),
    .O_1_0(n60_O_1_0),
    .O_1_1(n60_O_1_1),
    .O_1_2(n60_O_1_2),
    .O_2_0(n60_O_2_0),
    .O_2_1(n60_O_2_1),
    .O_2_2(n60_O_2_2),
    .O_3_0(n60_O_3_0),
    .O_3_1(n60_O_3_1),
    .O_3_2(n60_O_3_2),
    .O_4_0(n60_O_4_0),
    .O_4_1(n60_O_4_1),
    .O_4_2(n60_O_4_2),
    .O_5_0(n60_O_5_0),
    .O_5_1(n60_O_5_1),
    .O_5_2(n60_O_5_2),
    .O_6_0(n60_O_6_0),
    .O_6_1(n60_O_6_1),
    .O_6_2(n60_O_6_2),
    .O_7_0(n60_O_7_0),
    .O_7_1(n60_O_7_1),
    .O_7_2(n60_O_7_2),
    .O_8_0(n60_O_8_0),
    .O_8_1(n60_O_8_1),
    .O_8_2(n60_O_8_2),
    .O_9_0(n60_O_9_0),
    .O_9_1(n60_O_9_1),
    .O_9_2(n60_O_9_2),
    .O_10_0(n60_O_10_0),
    .O_10_1(n60_O_10_1),
    .O_10_2(n60_O_10_2),
    .O_11_0(n60_O_11_0),
    .O_11_1(n60_O_11_1),
    .O_11_2(n60_O_11_2),
    .O_12_0(n60_O_12_0),
    .O_12_1(n60_O_12_1),
    .O_12_2(n60_O_12_2),
    .O_13_0(n60_O_13_0),
    .O_13_1(n60_O_13_1),
    .O_13_2(n60_O_13_2),
    .O_14_0(n60_O_14_0),
    .O_14_1(n60_O_14_1),
    .O_14_2(n60_O_14_2),
    .O_15_0(n60_O_15_0),
    .O_15_1(n60_O_15_1),
    .O_15_2(n60_O_15_2)
  );
  Map2T_4 n61 ( // @[Top.scala 110:21]
    .valid_up(n61_valid_up),
    .valid_down(n61_valid_down),
    .I0_0_0(n61_I0_0_0),
    .I0_0_1(n61_I0_0_1),
    .I0_0_2(n61_I0_0_2),
    .I0_1_0(n61_I0_1_0),
    .I0_1_1(n61_I0_1_1),
    .I0_1_2(n61_I0_1_2),
    .I0_2_0(n61_I0_2_0),
    .I0_2_1(n61_I0_2_1),
    .I0_2_2(n61_I0_2_2),
    .I0_3_0(n61_I0_3_0),
    .I0_3_1(n61_I0_3_1),
    .I0_3_2(n61_I0_3_2),
    .I0_4_0(n61_I0_4_0),
    .I0_4_1(n61_I0_4_1),
    .I0_4_2(n61_I0_4_2),
    .I0_5_0(n61_I0_5_0),
    .I0_5_1(n61_I0_5_1),
    .I0_5_2(n61_I0_5_2),
    .I0_6_0(n61_I0_6_0),
    .I0_6_1(n61_I0_6_1),
    .I0_6_2(n61_I0_6_2),
    .I0_7_0(n61_I0_7_0),
    .I0_7_1(n61_I0_7_1),
    .I0_7_2(n61_I0_7_2),
    .I0_8_0(n61_I0_8_0),
    .I0_8_1(n61_I0_8_1),
    .I0_8_2(n61_I0_8_2),
    .I0_9_0(n61_I0_9_0),
    .I0_9_1(n61_I0_9_1),
    .I0_9_2(n61_I0_9_2),
    .I0_10_0(n61_I0_10_0),
    .I0_10_1(n61_I0_10_1),
    .I0_10_2(n61_I0_10_2),
    .I0_11_0(n61_I0_11_0),
    .I0_11_1(n61_I0_11_1),
    .I0_11_2(n61_I0_11_2),
    .I0_12_0(n61_I0_12_0),
    .I0_12_1(n61_I0_12_1),
    .I0_12_2(n61_I0_12_2),
    .I0_13_0(n61_I0_13_0),
    .I0_13_1(n61_I0_13_1),
    .I0_13_2(n61_I0_13_2),
    .I0_14_0(n61_I0_14_0),
    .I0_14_1(n61_I0_14_1),
    .I0_14_2(n61_I0_14_2),
    .I0_15_0(n61_I0_15_0),
    .I0_15_1(n61_I0_15_1),
    .I0_15_2(n61_I0_15_2),
    .I1_0_0(n61_I1_0_0),
    .I1_0_1(n61_I1_0_1),
    .I1_0_2(n61_I1_0_2),
    .I1_1_0(n61_I1_1_0),
    .I1_1_1(n61_I1_1_1),
    .I1_1_2(n61_I1_1_2),
    .I1_2_0(n61_I1_2_0),
    .I1_2_1(n61_I1_2_1),
    .I1_2_2(n61_I1_2_2),
    .I1_3_0(n61_I1_3_0),
    .I1_3_1(n61_I1_3_1),
    .I1_3_2(n61_I1_3_2),
    .I1_4_0(n61_I1_4_0),
    .I1_4_1(n61_I1_4_1),
    .I1_4_2(n61_I1_4_2),
    .I1_5_0(n61_I1_5_0),
    .I1_5_1(n61_I1_5_1),
    .I1_5_2(n61_I1_5_2),
    .I1_6_0(n61_I1_6_0),
    .I1_6_1(n61_I1_6_1),
    .I1_6_2(n61_I1_6_2),
    .I1_7_0(n61_I1_7_0),
    .I1_7_1(n61_I1_7_1),
    .I1_7_2(n61_I1_7_2),
    .I1_8_0(n61_I1_8_0),
    .I1_8_1(n61_I1_8_1),
    .I1_8_2(n61_I1_8_2),
    .I1_9_0(n61_I1_9_0),
    .I1_9_1(n61_I1_9_1),
    .I1_9_2(n61_I1_9_2),
    .I1_10_0(n61_I1_10_0),
    .I1_10_1(n61_I1_10_1),
    .I1_10_2(n61_I1_10_2),
    .I1_11_0(n61_I1_11_0),
    .I1_11_1(n61_I1_11_1),
    .I1_11_2(n61_I1_11_2),
    .I1_12_0(n61_I1_12_0),
    .I1_12_1(n61_I1_12_1),
    .I1_12_2(n61_I1_12_2),
    .I1_13_0(n61_I1_13_0),
    .I1_13_1(n61_I1_13_1),
    .I1_13_2(n61_I1_13_2),
    .I1_14_0(n61_I1_14_0),
    .I1_14_1(n61_I1_14_1),
    .I1_14_2(n61_I1_14_2),
    .I1_15_0(n61_I1_15_0),
    .I1_15_1(n61_I1_15_1),
    .I1_15_2(n61_I1_15_2),
    .O_0_0_0(n61_O_0_0_0),
    .O_0_0_1(n61_O_0_0_1),
    .O_0_0_2(n61_O_0_0_2),
    .O_0_1_0(n61_O_0_1_0),
    .O_0_1_1(n61_O_0_1_1),
    .O_0_1_2(n61_O_0_1_2),
    .O_1_0_0(n61_O_1_0_0),
    .O_1_0_1(n61_O_1_0_1),
    .O_1_0_2(n61_O_1_0_2),
    .O_1_1_0(n61_O_1_1_0),
    .O_1_1_1(n61_O_1_1_1),
    .O_1_1_2(n61_O_1_1_2),
    .O_2_0_0(n61_O_2_0_0),
    .O_2_0_1(n61_O_2_0_1),
    .O_2_0_2(n61_O_2_0_2),
    .O_2_1_0(n61_O_2_1_0),
    .O_2_1_1(n61_O_2_1_1),
    .O_2_1_2(n61_O_2_1_2),
    .O_3_0_0(n61_O_3_0_0),
    .O_3_0_1(n61_O_3_0_1),
    .O_3_0_2(n61_O_3_0_2),
    .O_3_1_0(n61_O_3_1_0),
    .O_3_1_1(n61_O_3_1_1),
    .O_3_1_2(n61_O_3_1_2),
    .O_4_0_0(n61_O_4_0_0),
    .O_4_0_1(n61_O_4_0_1),
    .O_4_0_2(n61_O_4_0_2),
    .O_4_1_0(n61_O_4_1_0),
    .O_4_1_1(n61_O_4_1_1),
    .O_4_1_2(n61_O_4_1_2),
    .O_5_0_0(n61_O_5_0_0),
    .O_5_0_1(n61_O_5_0_1),
    .O_5_0_2(n61_O_5_0_2),
    .O_5_1_0(n61_O_5_1_0),
    .O_5_1_1(n61_O_5_1_1),
    .O_5_1_2(n61_O_5_1_2),
    .O_6_0_0(n61_O_6_0_0),
    .O_6_0_1(n61_O_6_0_1),
    .O_6_0_2(n61_O_6_0_2),
    .O_6_1_0(n61_O_6_1_0),
    .O_6_1_1(n61_O_6_1_1),
    .O_6_1_2(n61_O_6_1_2),
    .O_7_0_0(n61_O_7_0_0),
    .O_7_0_1(n61_O_7_0_1),
    .O_7_0_2(n61_O_7_0_2),
    .O_7_1_0(n61_O_7_1_0),
    .O_7_1_1(n61_O_7_1_1),
    .O_7_1_2(n61_O_7_1_2),
    .O_8_0_0(n61_O_8_0_0),
    .O_8_0_1(n61_O_8_0_1),
    .O_8_0_2(n61_O_8_0_2),
    .O_8_1_0(n61_O_8_1_0),
    .O_8_1_1(n61_O_8_1_1),
    .O_8_1_2(n61_O_8_1_2),
    .O_9_0_0(n61_O_9_0_0),
    .O_9_0_1(n61_O_9_0_1),
    .O_9_0_2(n61_O_9_0_2),
    .O_9_1_0(n61_O_9_1_0),
    .O_9_1_1(n61_O_9_1_1),
    .O_9_1_2(n61_O_9_1_2),
    .O_10_0_0(n61_O_10_0_0),
    .O_10_0_1(n61_O_10_0_1),
    .O_10_0_2(n61_O_10_0_2),
    .O_10_1_0(n61_O_10_1_0),
    .O_10_1_1(n61_O_10_1_1),
    .O_10_1_2(n61_O_10_1_2),
    .O_11_0_0(n61_O_11_0_0),
    .O_11_0_1(n61_O_11_0_1),
    .O_11_0_2(n61_O_11_0_2),
    .O_11_1_0(n61_O_11_1_0),
    .O_11_1_1(n61_O_11_1_1),
    .O_11_1_2(n61_O_11_1_2),
    .O_12_0_0(n61_O_12_0_0),
    .O_12_0_1(n61_O_12_0_1),
    .O_12_0_2(n61_O_12_0_2),
    .O_12_1_0(n61_O_12_1_0),
    .O_12_1_1(n61_O_12_1_1),
    .O_12_1_2(n61_O_12_1_2),
    .O_13_0_0(n61_O_13_0_0),
    .O_13_0_1(n61_O_13_0_1),
    .O_13_0_2(n61_O_13_0_2),
    .O_13_1_0(n61_O_13_1_0),
    .O_13_1_1(n61_O_13_1_1),
    .O_13_1_2(n61_O_13_1_2),
    .O_14_0_0(n61_O_14_0_0),
    .O_14_0_1(n61_O_14_0_1),
    .O_14_0_2(n61_O_14_0_2),
    .O_14_1_0(n61_O_14_1_0),
    .O_14_1_1(n61_O_14_1_1),
    .O_14_1_2(n61_O_14_1_2),
    .O_15_0_0(n61_O_15_0_0),
    .O_15_0_1(n61_O_15_0_1),
    .O_15_0_2(n61_O_15_0_2),
    .O_15_1_0(n61_O_15_1_0),
    .O_15_1_1(n61_O_15_1_1),
    .O_15_1_2(n61_O_15_1_2)
  );
  ShiftTS_2 n68 ( // @[Top.scala 114:21]
    .clock(n68_clock),
    .reset(n68_reset),
    .valid_up(n68_valid_up),
    .valid_down(n68_valid_down),
    .I_0(n68_I_0),
    .I_1(n68_I_1),
    .I_2(n68_I_2),
    .I_3(n68_I_3),
    .I_4(n68_I_4),
    .I_5(n68_I_5),
    .I_6(n68_I_6),
    .I_7(n68_I_7),
    .I_8(n68_I_8),
    .I_9(n68_I_9),
    .I_10(n68_I_10),
    .I_11(n68_I_11),
    .I_12(n68_I_12),
    .I_13(n68_I_13),
    .I_14(n68_I_14),
    .I_15(n68_I_15),
    .O_0(n68_O_0),
    .O_1(n68_O_1),
    .O_2(n68_O_2),
    .O_3(n68_O_3),
    .O_4(n68_O_4),
    .O_5(n68_O_5),
    .O_6(n68_O_6),
    .O_7(n68_O_7),
    .O_8(n68_O_8),
    .O_9(n68_O_9),
    .O_10(n68_O_10),
    .O_11(n68_O_11),
    .O_12(n68_O_12),
    .O_13(n68_O_13),
    .O_14(n68_O_14),
    .O_15(n68_O_15)
  );
  ShiftTS_2 n69 ( // @[Top.scala 117:21]
    .clock(n69_clock),
    .reset(n69_reset),
    .valid_up(n69_valid_up),
    .valid_down(n69_valid_down),
    .I_0(n69_I_0),
    .I_1(n69_I_1),
    .I_2(n69_I_2),
    .I_3(n69_I_3),
    .I_4(n69_I_4),
    .I_5(n69_I_5),
    .I_6(n69_I_6),
    .I_7(n69_I_7),
    .I_8(n69_I_8),
    .I_9(n69_I_9),
    .I_10(n69_I_10),
    .I_11(n69_I_11),
    .I_12(n69_I_12),
    .I_13(n69_I_13),
    .I_14(n69_I_14),
    .I_15(n69_I_15),
    .O_0(n69_O_0),
    .O_1(n69_O_1),
    .O_2(n69_O_2),
    .O_3(n69_O_3),
    .O_4(n69_O_4),
    .O_5(n69_O_5),
    .O_6(n69_O_6),
    .O_7(n69_O_7),
    .O_8(n69_O_8),
    .O_9(n69_O_9),
    .O_10(n69_O_10),
    .O_11(n69_O_11),
    .O_12(n69_O_12),
    .O_13(n69_O_13),
    .O_14(n69_O_14),
    .O_15(n69_O_15)
  );
  FIFO n70 ( // @[Top.scala 120:21]
    .clock(n70_clock),
    .reset(n70_reset),
    .valid_up(n70_valid_up),
    .valid_down(n70_valid_down),
    .I_0(n70_I_0),
    .I_1(n70_I_1),
    .I_2(n70_I_2),
    .I_3(n70_I_3),
    .I_4(n70_I_4),
    .I_5(n70_I_5),
    .I_6(n70_I_6),
    .I_7(n70_I_7),
    .I_8(n70_I_8),
    .I_9(n70_I_9),
    .I_10(n70_I_10),
    .I_11(n70_I_11),
    .I_12(n70_I_12),
    .I_13(n70_I_13),
    .I_14(n70_I_14),
    .I_15(n70_I_15),
    .O_0(n70_O_0),
    .O_1(n70_O_1),
    .O_2(n70_O_2),
    .O_3(n70_O_3),
    .O_4(n70_O_4),
    .O_5(n70_O_5),
    .O_6(n70_O_6),
    .O_7(n70_O_7),
    .O_8(n70_O_8),
    .O_9(n70_O_9),
    .O_10(n70_O_10),
    .O_11(n70_O_11),
    .O_12(n70_O_12),
    .O_13(n70_O_13),
    .O_14(n70_O_14),
    .O_15(n70_O_15)
  );
  Map2T n71 ( // @[Top.scala 123:21]
    .valid_up(n71_valid_up),
    .valid_down(n71_valid_down),
    .I0_0(n71_I0_0),
    .I0_1(n71_I0_1),
    .I0_2(n71_I0_2),
    .I0_3(n71_I0_3),
    .I0_4(n71_I0_4),
    .I0_5(n71_I0_5),
    .I0_6(n71_I0_6),
    .I0_7(n71_I0_7),
    .I0_8(n71_I0_8),
    .I0_9(n71_I0_9),
    .I0_10(n71_I0_10),
    .I0_11(n71_I0_11),
    .I0_12(n71_I0_12),
    .I0_13(n71_I0_13),
    .I0_14(n71_I0_14),
    .I0_15(n71_I0_15),
    .I1_0(n71_I1_0),
    .I1_1(n71_I1_1),
    .I1_2(n71_I1_2),
    .I1_3(n71_I1_3),
    .I1_4(n71_I1_4),
    .I1_5(n71_I1_5),
    .I1_6(n71_I1_6),
    .I1_7(n71_I1_7),
    .I1_8(n71_I1_8),
    .I1_9(n71_I1_9),
    .I1_10(n71_I1_10),
    .I1_11(n71_I1_11),
    .I1_12(n71_I1_12),
    .I1_13(n71_I1_13),
    .I1_14(n71_I1_14),
    .I1_15(n71_I1_15),
    .O_0_0(n71_O_0_0),
    .O_0_1(n71_O_0_1),
    .O_1_0(n71_O_1_0),
    .O_1_1(n71_O_1_1),
    .O_2_0(n71_O_2_0),
    .O_2_1(n71_O_2_1),
    .O_3_0(n71_O_3_0),
    .O_3_1(n71_O_3_1),
    .O_4_0(n71_O_4_0),
    .O_4_1(n71_O_4_1),
    .O_5_0(n71_O_5_0),
    .O_5_1(n71_O_5_1),
    .O_6_0(n71_O_6_0),
    .O_6_1(n71_O_6_1),
    .O_7_0(n71_O_7_0),
    .O_7_1(n71_O_7_1),
    .O_8_0(n71_O_8_0),
    .O_8_1(n71_O_8_1),
    .O_9_0(n71_O_9_0),
    .O_9_1(n71_O_9_1),
    .O_10_0(n71_O_10_0),
    .O_10_1(n71_O_10_1),
    .O_11_0(n71_O_11_0),
    .O_11_1(n71_O_11_1),
    .O_12_0(n71_O_12_0),
    .O_12_1(n71_O_12_1),
    .O_13_0(n71_O_13_0),
    .O_13_1(n71_O_13_1),
    .O_14_0(n71_O_14_0),
    .O_14_1(n71_O_14_1),
    .O_15_0(n71_O_15_0),
    .O_15_1(n71_O_15_1)
  );
  FIFO_2 n78 ( // @[Top.scala 127:21]
    .clock(n78_clock),
    .reset(n78_reset),
    .valid_up(n78_valid_up),
    .valid_down(n78_valid_down),
    .I_0(n78_I_0),
    .I_1(n78_I_1),
    .I_2(n78_I_2),
    .I_3(n78_I_3),
    .I_4(n78_I_4),
    .I_5(n78_I_5),
    .I_6(n78_I_6),
    .I_7(n78_I_7),
    .I_8(n78_I_8),
    .I_9(n78_I_9),
    .I_10(n78_I_10),
    .I_11(n78_I_11),
    .I_12(n78_I_12),
    .I_13(n78_I_13),
    .I_14(n78_I_14),
    .I_15(n78_I_15),
    .O_0(n78_O_0),
    .O_1(n78_O_1),
    .O_2(n78_O_2),
    .O_3(n78_O_3),
    .O_4(n78_O_4),
    .O_5(n78_O_5),
    .O_6(n78_O_6),
    .O_7(n78_O_7),
    .O_8(n78_O_8),
    .O_9(n78_O_9),
    .O_10(n78_O_10),
    .O_11(n78_O_11),
    .O_12(n78_O_12),
    .O_13(n78_O_13),
    .O_14(n78_O_14),
    .O_15(n78_O_15)
  );
  Map2T_1 n79 ( // @[Top.scala 130:21]
    .valid_up(n79_valid_up),
    .valid_down(n79_valid_down),
    .I0_0_0(n79_I0_0_0),
    .I0_0_1(n79_I0_0_1),
    .I0_1_0(n79_I0_1_0),
    .I0_1_1(n79_I0_1_1),
    .I0_2_0(n79_I0_2_0),
    .I0_2_1(n79_I0_2_1),
    .I0_3_0(n79_I0_3_0),
    .I0_3_1(n79_I0_3_1),
    .I0_4_0(n79_I0_4_0),
    .I0_4_1(n79_I0_4_1),
    .I0_5_0(n79_I0_5_0),
    .I0_5_1(n79_I0_5_1),
    .I0_6_0(n79_I0_6_0),
    .I0_6_1(n79_I0_6_1),
    .I0_7_0(n79_I0_7_0),
    .I0_7_1(n79_I0_7_1),
    .I0_8_0(n79_I0_8_0),
    .I0_8_1(n79_I0_8_1),
    .I0_9_0(n79_I0_9_0),
    .I0_9_1(n79_I0_9_1),
    .I0_10_0(n79_I0_10_0),
    .I0_10_1(n79_I0_10_1),
    .I0_11_0(n79_I0_11_0),
    .I0_11_1(n79_I0_11_1),
    .I0_12_0(n79_I0_12_0),
    .I0_12_1(n79_I0_12_1),
    .I0_13_0(n79_I0_13_0),
    .I0_13_1(n79_I0_13_1),
    .I0_14_0(n79_I0_14_0),
    .I0_14_1(n79_I0_14_1),
    .I0_15_0(n79_I0_15_0),
    .I0_15_1(n79_I0_15_1),
    .I1_0(n79_I1_0),
    .I1_1(n79_I1_1),
    .I1_2(n79_I1_2),
    .I1_3(n79_I1_3),
    .I1_4(n79_I1_4),
    .I1_5(n79_I1_5),
    .I1_6(n79_I1_6),
    .I1_7(n79_I1_7),
    .I1_8(n79_I1_8),
    .I1_9(n79_I1_9),
    .I1_10(n79_I1_10),
    .I1_11(n79_I1_11),
    .I1_12(n79_I1_12),
    .I1_13(n79_I1_13),
    .I1_14(n79_I1_14),
    .I1_15(n79_I1_15),
    .O_0_0(n79_O_0_0),
    .O_0_1(n79_O_0_1),
    .O_0_2(n79_O_0_2),
    .O_1_0(n79_O_1_0),
    .O_1_1(n79_O_1_1),
    .O_1_2(n79_O_1_2),
    .O_2_0(n79_O_2_0),
    .O_2_1(n79_O_2_1),
    .O_2_2(n79_O_2_2),
    .O_3_0(n79_O_3_0),
    .O_3_1(n79_O_3_1),
    .O_3_2(n79_O_3_2),
    .O_4_0(n79_O_4_0),
    .O_4_1(n79_O_4_1),
    .O_4_2(n79_O_4_2),
    .O_5_0(n79_O_5_0),
    .O_5_1(n79_O_5_1),
    .O_5_2(n79_O_5_2),
    .O_6_0(n79_O_6_0),
    .O_6_1(n79_O_6_1),
    .O_6_2(n79_O_6_2),
    .O_7_0(n79_O_7_0),
    .O_7_1(n79_O_7_1),
    .O_7_2(n79_O_7_2),
    .O_8_0(n79_O_8_0),
    .O_8_1(n79_O_8_1),
    .O_8_2(n79_O_8_2),
    .O_9_0(n79_O_9_0),
    .O_9_1(n79_O_9_1),
    .O_9_2(n79_O_9_2),
    .O_10_0(n79_O_10_0),
    .O_10_1(n79_O_10_1),
    .O_10_2(n79_O_10_2),
    .O_11_0(n79_O_11_0),
    .O_11_1(n79_O_11_1),
    .O_11_2(n79_O_11_2),
    .O_12_0(n79_O_12_0),
    .O_12_1(n79_O_12_1),
    .O_12_2(n79_O_12_2),
    .O_13_0(n79_O_13_0),
    .O_13_1(n79_O_13_1),
    .O_13_2(n79_O_13_2),
    .O_14_0(n79_O_14_0),
    .O_14_1(n79_O_14_1),
    .O_14_2(n79_O_14_2),
    .O_15_0(n79_O_15_0),
    .O_15_1(n79_O_15_1),
    .O_15_2(n79_O_15_2)
  );
  MapT n88 ( // @[Top.scala 134:21]
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0(n88_I_0_0),
    .I_0_1(n88_I_0_1),
    .I_0_2(n88_I_0_2),
    .I_1_0(n88_I_1_0),
    .I_1_1(n88_I_1_1),
    .I_1_2(n88_I_1_2),
    .I_2_0(n88_I_2_0),
    .I_2_1(n88_I_2_1),
    .I_2_2(n88_I_2_2),
    .I_3_0(n88_I_3_0),
    .I_3_1(n88_I_3_1),
    .I_3_2(n88_I_3_2),
    .I_4_0(n88_I_4_0),
    .I_4_1(n88_I_4_1),
    .I_4_2(n88_I_4_2),
    .I_5_0(n88_I_5_0),
    .I_5_1(n88_I_5_1),
    .I_5_2(n88_I_5_2),
    .I_6_0(n88_I_6_0),
    .I_6_1(n88_I_6_1),
    .I_6_2(n88_I_6_2),
    .I_7_0(n88_I_7_0),
    .I_7_1(n88_I_7_1),
    .I_7_2(n88_I_7_2),
    .I_8_0(n88_I_8_0),
    .I_8_1(n88_I_8_1),
    .I_8_2(n88_I_8_2),
    .I_9_0(n88_I_9_0),
    .I_9_1(n88_I_9_1),
    .I_9_2(n88_I_9_2),
    .I_10_0(n88_I_10_0),
    .I_10_1(n88_I_10_1),
    .I_10_2(n88_I_10_2),
    .I_11_0(n88_I_11_0),
    .I_11_1(n88_I_11_1),
    .I_11_2(n88_I_11_2),
    .I_12_0(n88_I_12_0),
    .I_12_1(n88_I_12_1),
    .I_12_2(n88_I_12_2),
    .I_13_0(n88_I_13_0),
    .I_13_1(n88_I_13_1),
    .I_13_2(n88_I_13_2),
    .I_14_0(n88_I_14_0),
    .I_14_1(n88_I_14_1),
    .I_14_2(n88_I_14_2),
    .I_15_0(n88_I_15_0),
    .I_15_1(n88_I_15_1),
    .I_15_2(n88_I_15_2),
    .O_0_0_0(n88_O_0_0_0),
    .O_0_0_1(n88_O_0_0_1),
    .O_0_0_2(n88_O_0_0_2),
    .O_1_0_0(n88_O_1_0_0),
    .O_1_0_1(n88_O_1_0_1),
    .O_1_0_2(n88_O_1_0_2),
    .O_2_0_0(n88_O_2_0_0),
    .O_2_0_1(n88_O_2_0_1),
    .O_2_0_2(n88_O_2_0_2),
    .O_3_0_0(n88_O_3_0_0),
    .O_3_0_1(n88_O_3_0_1),
    .O_3_0_2(n88_O_3_0_2),
    .O_4_0_0(n88_O_4_0_0),
    .O_4_0_1(n88_O_4_0_1),
    .O_4_0_2(n88_O_4_0_2),
    .O_5_0_0(n88_O_5_0_0),
    .O_5_0_1(n88_O_5_0_1),
    .O_5_0_2(n88_O_5_0_2),
    .O_6_0_0(n88_O_6_0_0),
    .O_6_0_1(n88_O_6_0_1),
    .O_6_0_2(n88_O_6_0_2),
    .O_7_0_0(n88_O_7_0_0),
    .O_7_0_1(n88_O_7_0_1),
    .O_7_0_2(n88_O_7_0_2),
    .O_8_0_0(n88_O_8_0_0),
    .O_8_0_1(n88_O_8_0_1),
    .O_8_0_2(n88_O_8_0_2),
    .O_9_0_0(n88_O_9_0_0),
    .O_9_0_1(n88_O_9_0_1),
    .O_9_0_2(n88_O_9_0_2),
    .O_10_0_0(n88_O_10_0_0),
    .O_10_0_1(n88_O_10_0_1),
    .O_10_0_2(n88_O_10_0_2),
    .O_11_0_0(n88_O_11_0_0),
    .O_11_0_1(n88_O_11_0_1),
    .O_11_0_2(n88_O_11_0_2),
    .O_12_0_0(n88_O_12_0_0),
    .O_12_0_1(n88_O_12_0_1),
    .O_12_0_2(n88_O_12_0_2),
    .O_13_0_0(n88_O_13_0_0),
    .O_13_0_1(n88_O_13_0_1),
    .O_13_0_2(n88_O_13_0_2),
    .O_14_0_0(n88_O_14_0_0),
    .O_14_0_1(n88_O_14_0_1),
    .O_14_0_2(n88_O_14_0_2),
    .O_15_0_0(n88_O_15_0_0),
    .O_15_0_1(n88_O_15_0_1),
    .O_15_0_2(n88_O_15_0_2)
  );
  MapT_1 n95 ( // @[Top.scala 137:21]
    .valid_up(n95_valid_up),
    .valid_down(n95_valid_down),
    .I_0_0_0(n95_I_0_0_0),
    .I_0_0_1(n95_I_0_0_1),
    .I_0_0_2(n95_I_0_0_2),
    .I_1_0_0(n95_I_1_0_0),
    .I_1_0_1(n95_I_1_0_1),
    .I_1_0_2(n95_I_1_0_2),
    .I_2_0_0(n95_I_2_0_0),
    .I_2_0_1(n95_I_2_0_1),
    .I_2_0_2(n95_I_2_0_2),
    .I_3_0_0(n95_I_3_0_0),
    .I_3_0_1(n95_I_3_0_1),
    .I_3_0_2(n95_I_3_0_2),
    .I_4_0_0(n95_I_4_0_0),
    .I_4_0_1(n95_I_4_0_1),
    .I_4_0_2(n95_I_4_0_2),
    .I_5_0_0(n95_I_5_0_0),
    .I_5_0_1(n95_I_5_0_1),
    .I_5_0_2(n95_I_5_0_2),
    .I_6_0_0(n95_I_6_0_0),
    .I_6_0_1(n95_I_6_0_1),
    .I_6_0_2(n95_I_6_0_2),
    .I_7_0_0(n95_I_7_0_0),
    .I_7_0_1(n95_I_7_0_1),
    .I_7_0_2(n95_I_7_0_2),
    .I_8_0_0(n95_I_8_0_0),
    .I_8_0_1(n95_I_8_0_1),
    .I_8_0_2(n95_I_8_0_2),
    .I_9_0_0(n95_I_9_0_0),
    .I_9_0_1(n95_I_9_0_1),
    .I_9_0_2(n95_I_9_0_2),
    .I_10_0_0(n95_I_10_0_0),
    .I_10_0_1(n95_I_10_0_1),
    .I_10_0_2(n95_I_10_0_2),
    .I_11_0_0(n95_I_11_0_0),
    .I_11_0_1(n95_I_11_0_1),
    .I_11_0_2(n95_I_11_0_2),
    .I_12_0_0(n95_I_12_0_0),
    .I_12_0_1(n95_I_12_0_1),
    .I_12_0_2(n95_I_12_0_2),
    .I_13_0_0(n95_I_13_0_0),
    .I_13_0_1(n95_I_13_0_1),
    .I_13_0_2(n95_I_13_0_2),
    .I_14_0_0(n95_I_14_0_0),
    .I_14_0_1(n95_I_14_0_1),
    .I_14_0_2(n95_I_14_0_2),
    .I_15_0_0(n95_I_15_0_0),
    .I_15_0_1(n95_I_15_0_1),
    .I_15_0_2(n95_I_15_0_2),
    .O_0_0(n95_O_0_0),
    .O_0_1(n95_O_0_1),
    .O_0_2(n95_O_0_2),
    .O_1_0(n95_O_1_0),
    .O_1_1(n95_O_1_1),
    .O_1_2(n95_O_1_2),
    .O_2_0(n95_O_2_0),
    .O_2_1(n95_O_2_1),
    .O_2_2(n95_O_2_2),
    .O_3_0(n95_O_3_0),
    .O_3_1(n95_O_3_1),
    .O_3_2(n95_O_3_2),
    .O_4_0(n95_O_4_0),
    .O_4_1(n95_O_4_1),
    .O_4_2(n95_O_4_2),
    .O_5_0(n95_O_5_0),
    .O_5_1(n95_O_5_1),
    .O_5_2(n95_O_5_2),
    .O_6_0(n95_O_6_0),
    .O_6_1(n95_O_6_1),
    .O_6_2(n95_O_6_2),
    .O_7_0(n95_O_7_0),
    .O_7_1(n95_O_7_1),
    .O_7_2(n95_O_7_2),
    .O_8_0(n95_O_8_0),
    .O_8_1(n95_O_8_1),
    .O_8_2(n95_O_8_2),
    .O_9_0(n95_O_9_0),
    .O_9_1(n95_O_9_1),
    .O_9_2(n95_O_9_2),
    .O_10_0(n95_O_10_0),
    .O_10_1(n95_O_10_1),
    .O_10_2(n95_O_10_2),
    .O_11_0(n95_O_11_0),
    .O_11_1(n95_O_11_1),
    .O_11_2(n95_O_11_2),
    .O_12_0(n95_O_12_0),
    .O_12_1(n95_O_12_1),
    .O_12_2(n95_O_12_2),
    .O_13_0(n95_O_13_0),
    .O_13_1(n95_O_13_1),
    .O_13_2(n95_O_13_2),
    .O_14_0(n95_O_14_0),
    .O_14_1(n95_O_14_1),
    .O_14_2(n95_O_14_2),
    .O_15_0(n95_O_15_0),
    .O_15_1(n95_O_15_1),
    .O_15_2(n95_O_15_2)
  );
  FIFO_8 n96 ( // @[Top.scala 140:21]
    .clock(n96_clock),
    .reset(n96_reset),
    .valid_up(n96_valid_up),
    .valid_down(n96_valid_down),
    .I_0_0(n96_I_0_0),
    .I_0_1(n96_I_0_1),
    .I_0_2(n96_I_0_2),
    .I_1_0(n96_I_1_0),
    .I_1_1(n96_I_1_1),
    .I_1_2(n96_I_1_2),
    .I_2_0(n96_I_2_0),
    .I_2_1(n96_I_2_1),
    .I_2_2(n96_I_2_2),
    .I_3_0(n96_I_3_0),
    .I_3_1(n96_I_3_1),
    .I_3_2(n96_I_3_2),
    .I_4_0(n96_I_4_0),
    .I_4_1(n96_I_4_1),
    .I_4_2(n96_I_4_2),
    .I_5_0(n96_I_5_0),
    .I_5_1(n96_I_5_1),
    .I_5_2(n96_I_5_2),
    .I_6_0(n96_I_6_0),
    .I_6_1(n96_I_6_1),
    .I_6_2(n96_I_6_2),
    .I_7_0(n96_I_7_0),
    .I_7_1(n96_I_7_1),
    .I_7_2(n96_I_7_2),
    .I_8_0(n96_I_8_0),
    .I_8_1(n96_I_8_1),
    .I_8_2(n96_I_8_2),
    .I_9_0(n96_I_9_0),
    .I_9_1(n96_I_9_1),
    .I_9_2(n96_I_9_2),
    .I_10_0(n96_I_10_0),
    .I_10_1(n96_I_10_1),
    .I_10_2(n96_I_10_2),
    .I_11_0(n96_I_11_0),
    .I_11_1(n96_I_11_1),
    .I_11_2(n96_I_11_2),
    .I_12_0(n96_I_12_0),
    .I_12_1(n96_I_12_1),
    .I_12_2(n96_I_12_2),
    .I_13_0(n96_I_13_0),
    .I_13_1(n96_I_13_1),
    .I_13_2(n96_I_13_2),
    .I_14_0(n96_I_14_0),
    .I_14_1(n96_I_14_1),
    .I_14_2(n96_I_14_2),
    .I_15_0(n96_I_15_0),
    .I_15_1(n96_I_15_1),
    .I_15_2(n96_I_15_2),
    .O_0_0(n96_O_0_0),
    .O_0_1(n96_O_0_1),
    .O_0_2(n96_O_0_2),
    .O_1_0(n96_O_1_0),
    .O_1_1(n96_O_1_1),
    .O_1_2(n96_O_1_2),
    .O_2_0(n96_O_2_0),
    .O_2_1(n96_O_2_1),
    .O_2_2(n96_O_2_2),
    .O_3_0(n96_O_3_0),
    .O_3_1(n96_O_3_1),
    .O_3_2(n96_O_3_2),
    .O_4_0(n96_O_4_0),
    .O_4_1(n96_O_4_1),
    .O_4_2(n96_O_4_2),
    .O_5_0(n96_O_5_0),
    .O_5_1(n96_O_5_1),
    .O_5_2(n96_O_5_2),
    .O_6_0(n96_O_6_0),
    .O_6_1(n96_O_6_1),
    .O_6_2(n96_O_6_2),
    .O_7_0(n96_O_7_0),
    .O_7_1(n96_O_7_1),
    .O_7_2(n96_O_7_2),
    .O_8_0(n96_O_8_0),
    .O_8_1(n96_O_8_1),
    .O_8_2(n96_O_8_2),
    .O_9_0(n96_O_9_0),
    .O_9_1(n96_O_9_1),
    .O_9_2(n96_O_9_2),
    .O_10_0(n96_O_10_0),
    .O_10_1(n96_O_10_1),
    .O_10_2(n96_O_10_2),
    .O_11_0(n96_O_11_0),
    .O_11_1(n96_O_11_1),
    .O_11_2(n96_O_11_2),
    .O_12_0(n96_O_12_0),
    .O_12_1(n96_O_12_1),
    .O_12_2(n96_O_12_2),
    .O_13_0(n96_O_13_0),
    .O_13_1(n96_O_13_1),
    .O_13_2(n96_O_13_2),
    .O_14_0(n96_O_14_0),
    .O_14_1(n96_O_14_1),
    .O_14_2(n96_O_14_2),
    .O_15_0(n96_O_15_0),
    .O_15_1(n96_O_15_1),
    .O_15_2(n96_O_15_2)
  );
  Map2T_7 n97 ( // @[Top.scala 143:21]
    .valid_up(n97_valid_up),
    .valid_down(n97_valid_down),
    .I0_0_0_0(n97_I0_0_0_0),
    .I0_0_0_1(n97_I0_0_0_1),
    .I0_0_0_2(n97_I0_0_0_2),
    .I0_0_1_0(n97_I0_0_1_0),
    .I0_0_1_1(n97_I0_0_1_1),
    .I0_0_1_2(n97_I0_0_1_2),
    .I0_1_0_0(n97_I0_1_0_0),
    .I0_1_0_1(n97_I0_1_0_1),
    .I0_1_0_2(n97_I0_1_0_2),
    .I0_1_1_0(n97_I0_1_1_0),
    .I0_1_1_1(n97_I0_1_1_1),
    .I0_1_1_2(n97_I0_1_1_2),
    .I0_2_0_0(n97_I0_2_0_0),
    .I0_2_0_1(n97_I0_2_0_1),
    .I0_2_0_2(n97_I0_2_0_2),
    .I0_2_1_0(n97_I0_2_1_0),
    .I0_2_1_1(n97_I0_2_1_1),
    .I0_2_1_2(n97_I0_2_1_2),
    .I0_3_0_0(n97_I0_3_0_0),
    .I0_3_0_1(n97_I0_3_0_1),
    .I0_3_0_2(n97_I0_3_0_2),
    .I0_3_1_0(n97_I0_3_1_0),
    .I0_3_1_1(n97_I0_3_1_1),
    .I0_3_1_2(n97_I0_3_1_2),
    .I0_4_0_0(n97_I0_4_0_0),
    .I0_4_0_1(n97_I0_4_0_1),
    .I0_4_0_2(n97_I0_4_0_2),
    .I0_4_1_0(n97_I0_4_1_0),
    .I0_4_1_1(n97_I0_4_1_1),
    .I0_4_1_2(n97_I0_4_1_2),
    .I0_5_0_0(n97_I0_5_0_0),
    .I0_5_0_1(n97_I0_5_0_1),
    .I0_5_0_2(n97_I0_5_0_2),
    .I0_5_1_0(n97_I0_5_1_0),
    .I0_5_1_1(n97_I0_5_1_1),
    .I0_5_1_2(n97_I0_5_1_2),
    .I0_6_0_0(n97_I0_6_0_0),
    .I0_6_0_1(n97_I0_6_0_1),
    .I0_6_0_2(n97_I0_6_0_2),
    .I0_6_1_0(n97_I0_6_1_0),
    .I0_6_1_1(n97_I0_6_1_1),
    .I0_6_1_2(n97_I0_6_1_2),
    .I0_7_0_0(n97_I0_7_0_0),
    .I0_7_0_1(n97_I0_7_0_1),
    .I0_7_0_2(n97_I0_7_0_2),
    .I0_7_1_0(n97_I0_7_1_0),
    .I0_7_1_1(n97_I0_7_1_1),
    .I0_7_1_2(n97_I0_7_1_2),
    .I0_8_0_0(n97_I0_8_0_0),
    .I0_8_0_1(n97_I0_8_0_1),
    .I0_8_0_2(n97_I0_8_0_2),
    .I0_8_1_0(n97_I0_8_1_0),
    .I0_8_1_1(n97_I0_8_1_1),
    .I0_8_1_2(n97_I0_8_1_2),
    .I0_9_0_0(n97_I0_9_0_0),
    .I0_9_0_1(n97_I0_9_0_1),
    .I0_9_0_2(n97_I0_9_0_2),
    .I0_9_1_0(n97_I0_9_1_0),
    .I0_9_1_1(n97_I0_9_1_1),
    .I0_9_1_2(n97_I0_9_1_2),
    .I0_10_0_0(n97_I0_10_0_0),
    .I0_10_0_1(n97_I0_10_0_1),
    .I0_10_0_2(n97_I0_10_0_2),
    .I0_10_1_0(n97_I0_10_1_0),
    .I0_10_1_1(n97_I0_10_1_1),
    .I0_10_1_2(n97_I0_10_1_2),
    .I0_11_0_0(n97_I0_11_0_0),
    .I0_11_0_1(n97_I0_11_0_1),
    .I0_11_0_2(n97_I0_11_0_2),
    .I0_11_1_0(n97_I0_11_1_0),
    .I0_11_1_1(n97_I0_11_1_1),
    .I0_11_1_2(n97_I0_11_1_2),
    .I0_12_0_0(n97_I0_12_0_0),
    .I0_12_0_1(n97_I0_12_0_1),
    .I0_12_0_2(n97_I0_12_0_2),
    .I0_12_1_0(n97_I0_12_1_0),
    .I0_12_1_1(n97_I0_12_1_1),
    .I0_12_1_2(n97_I0_12_1_2),
    .I0_13_0_0(n97_I0_13_0_0),
    .I0_13_0_1(n97_I0_13_0_1),
    .I0_13_0_2(n97_I0_13_0_2),
    .I0_13_1_0(n97_I0_13_1_0),
    .I0_13_1_1(n97_I0_13_1_1),
    .I0_13_1_2(n97_I0_13_1_2),
    .I0_14_0_0(n97_I0_14_0_0),
    .I0_14_0_1(n97_I0_14_0_1),
    .I0_14_0_2(n97_I0_14_0_2),
    .I0_14_1_0(n97_I0_14_1_0),
    .I0_14_1_1(n97_I0_14_1_1),
    .I0_14_1_2(n97_I0_14_1_2),
    .I0_15_0_0(n97_I0_15_0_0),
    .I0_15_0_1(n97_I0_15_0_1),
    .I0_15_0_2(n97_I0_15_0_2),
    .I0_15_1_0(n97_I0_15_1_0),
    .I0_15_1_1(n97_I0_15_1_1),
    .I0_15_1_2(n97_I0_15_1_2),
    .I1_0_0(n97_I1_0_0),
    .I1_0_1(n97_I1_0_1),
    .I1_0_2(n97_I1_0_2),
    .I1_1_0(n97_I1_1_0),
    .I1_1_1(n97_I1_1_1),
    .I1_1_2(n97_I1_1_2),
    .I1_2_0(n97_I1_2_0),
    .I1_2_1(n97_I1_2_1),
    .I1_2_2(n97_I1_2_2),
    .I1_3_0(n97_I1_3_0),
    .I1_3_1(n97_I1_3_1),
    .I1_3_2(n97_I1_3_2),
    .I1_4_0(n97_I1_4_0),
    .I1_4_1(n97_I1_4_1),
    .I1_4_2(n97_I1_4_2),
    .I1_5_0(n97_I1_5_0),
    .I1_5_1(n97_I1_5_1),
    .I1_5_2(n97_I1_5_2),
    .I1_6_0(n97_I1_6_0),
    .I1_6_1(n97_I1_6_1),
    .I1_6_2(n97_I1_6_2),
    .I1_7_0(n97_I1_7_0),
    .I1_7_1(n97_I1_7_1),
    .I1_7_2(n97_I1_7_2),
    .I1_8_0(n97_I1_8_0),
    .I1_8_1(n97_I1_8_1),
    .I1_8_2(n97_I1_8_2),
    .I1_9_0(n97_I1_9_0),
    .I1_9_1(n97_I1_9_1),
    .I1_9_2(n97_I1_9_2),
    .I1_10_0(n97_I1_10_0),
    .I1_10_1(n97_I1_10_1),
    .I1_10_2(n97_I1_10_2),
    .I1_11_0(n97_I1_11_0),
    .I1_11_1(n97_I1_11_1),
    .I1_11_2(n97_I1_11_2),
    .I1_12_0(n97_I1_12_0),
    .I1_12_1(n97_I1_12_1),
    .I1_12_2(n97_I1_12_2),
    .I1_13_0(n97_I1_13_0),
    .I1_13_1(n97_I1_13_1),
    .I1_13_2(n97_I1_13_2),
    .I1_14_0(n97_I1_14_0),
    .I1_14_1(n97_I1_14_1),
    .I1_14_2(n97_I1_14_2),
    .I1_15_0(n97_I1_15_0),
    .I1_15_1(n97_I1_15_1),
    .I1_15_2(n97_I1_15_2),
    .O_0_0_0(n97_O_0_0_0),
    .O_0_0_1(n97_O_0_0_1),
    .O_0_0_2(n97_O_0_0_2),
    .O_0_1_0(n97_O_0_1_0),
    .O_0_1_1(n97_O_0_1_1),
    .O_0_1_2(n97_O_0_1_2),
    .O_0_2_0(n97_O_0_2_0),
    .O_0_2_1(n97_O_0_2_1),
    .O_0_2_2(n97_O_0_2_2),
    .O_1_0_0(n97_O_1_0_0),
    .O_1_0_1(n97_O_1_0_1),
    .O_1_0_2(n97_O_1_0_2),
    .O_1_1_0(n97_O_1_1_0),
    .O_1_1_1(n97_O_1_1_1),
    .O_1_1_2(n97_O_1_1_2),
    .O_1_2_0(n97_O_1_2_0),
    .O_1_2_1(n97_O_1_2_1),
    .O_1_2_2(n97_O_1_2_2),
    .O_2_0_0(n97_O_2_0_0),
    .O_2_0_1(n97_O_2_0_1),
    .O_2_0_2(n97_O_2_0_2),
    .O_2_1_0(n97_O_2_1_0),
    .O_2_1_1(n97_O_2_1_1),
    .O_2_1_2(n97_O_2_1_2),
    .O_2_2_0(n97_O_2_2_0),
    .O_2_2_1(n97_O_2_2_1),
    .O_2_2_2(n97_O_2_2_2),
    .O_3_0_0(n97_O_3_0_0),
    .O_3_0_1(n97_O_3_0_1),
    .O_3_0_2(n97_O_3_0_2),
    .O_3_1_0(n97_O_3_1_0),
    .O_3_1_1(n97_O_3_1_1),
    .O_3_1_2(n97_O_3_1_2),
    .O_3_2_0(n97_O_3_2_0),
    .O_3_2_1(n97_O_3_2_1),
    .O_3_2_2(n97_O_3_2_2),
    .O_4_0_0(n97_O_4_0_0),
    .O_4_0_1(n97_O_4_0_1),
    .O_4_0_2(n97_O_4_0_2),
    .O_4_1_0(n97_O_4_1_0),
    .O_4_1_1(n97_O_4_1_1),
    .O_4_1_2(n97_O_4_1_2),
    .O_4_2_0(n97_O_4_2_0),
    .O_4_2_1(n97_O_4_2_1),
    .O_4_2_2(n97_O_4_2_2),
    .O_5_0_0(n97_O_5_0_0),
    .O_5_0_1(n97_O_5_0_1),
    .O_5_0_2(n97_O_5_0_2),
    .O_5_1_0(n97_O_5_1_0),
    .O_5_1_1(n97_O_5_1_1),
    .O_5_1_2(n97_O_5_1_2),
    .O_5_2_0(n97_O_5_2_0),
    .O_5_2_1(n97_O_5_2_1),
    .O_5_2_2(n97_O_5_2_2),
    .O_6_0_0(n97_O_6_0_0),
    .O_6_0_1(n97_O_6_0_1),
    .O_6_0_2(n97_O_6_0_2),
    .O_6_1_0(n97_O_6_1_0),
    .O_6_1_1(n97_O_6_1_1),
    .O_6_1_2(n97_O_6_1_2),
    .O_6_2_0(n97_O_6_2_0),
    .O_6_2_1(n97_O_6_2_1),
    .O_6_2_2(n97_O_6_2_2),
    .O_7_0_0(n97_O_7_0_0),
    .O_7_0_1(n97_O_7_0_1),
    .O_7_0_2(n97_O_7_0_2),
    .O_7_1_0(n97_O_7_1_0),
    .O_7_1_1(n97_O_7_1_1),
    .O_7_1_2(n97_O_7_1_2),
    .O_7_2_0(n97_O_7_2_0),
    .O_7_2_1(n97_O_7_2_1),
    .O_7_2_2(n97_O_7_2_2),
    .O_8_0_0(n97_O_8_0_0),
    .O_8_0_1(n97_O_8_0_1),
    .O_8_0_2(n97_O_8_0_2),
    .O_8_1_0(n97_O_8_1_0),
    .O_8_1_1(n97_O_8_1_1),
    .O_8_1_2(n97_O_8_1_2),
    .O_8_2_0(n97_O_8_2_0),
    .O_8_2_1(n97_O_8_2_1),
    .O_8_2_2(n97_O_8_2_2),
    .O_9_0_0(n97_O_9_0_0),
    .O_9_0_1(n97_O_9_0_1),
    .O_9_0_2(n97_O_9_0_2),
    .O_9_1_0(n97_O_9_1_0),
    .O_9_1_1(n97_O_9_1_1),
    .O_9_1_2(n97_O_9_1_2),
    .O_9_2_0(n97_O_9_2_0),
    .O_9_2_1(n97_O_9_2_1),
    .O_9_2_2(n97_O_9_2_2),
    .O_10_0_0(n97_O_10_0_0),
    .O_10_0_1(n97_O_10_0_1),
    .O_10_0_2(n97_O_10_0_2),
    .O_10_1_0(n97_O_10_1_0),
    .O_10_1_1(n97_O_10_1_1),
    .O_10_1_2(n97_O_10_1_2),
    .O_10_2_0(n97_O_10_2_0),
    .O_10_2_1(n97_O_10_2_1),
    .O_10_2_2(n97_O_10_2_2),
    .O_11_0_0(n97_O_11_0_0),
    .O_11_0_1(n97_O_11_0_1),
    .O_11_0_2(n97_O_11_0_2),
    .O_11_1_0(n97_O_11_1_0),
    .O_11_1_1(n97_O_11_1_1),
    .O_11_1_2(n97_O_11_1_2),
    .O_11_2_0(n97_O_11_2_0),
    .O_11_2_1(n97_O_11_2_1),
    .O_11_2_2(n97_O_11_2_2),
    .O_12_0_0(n97_O_12_0_0),
    .O_12_0_1(n97_O_12_0_1),
    .O_12_0_2(n97_O_12_0_2),
    .O_12_1_0(n97_O_12_1_0),
    .O_12_1_1(n97_O_12_1_1),
    .O_12_1_2(n97_O_12_1_2),
    .O_12_2_0(n97_O_12_2_0),
    .O_12_2_1(n97_O_12_2_1),
    .O_12_2_2(n97_O_12_2_2),
    .O_13_0_0(n97_O_13_0_0),
    .O_13_0_1(n97_O_13_0_1),
    .O_13_0_2(n97_O_13_0_2),
    .O_13_1_0(n97_O_13_1_0),
    .O_13_1_1(n97_O_13_1_1),
    .O_13_1_2(n97_O_13_1_2),
    .O_13_2_0(n97_O_13_2_0),
    .O_13_2_1(n97_O_13_2_1),
    .O_13_2_2(n97_O_13_2_2),
    .O_14_0_0(n97_O_14_0_0),
    .O_14_0_1(n97_O_14_0_1),
    .O_14_0_2(n97_O_14_0_2),
    .O_14_1_0(n97_O_14_1_0),
    .O_14_1_1(n97_O_14_1_1),
    .O_14_1_2(n97_O_14_1_2),
    .O_14_2_0(n97_O_14_2_0),
    .O_14_2_1(n97_O_14_2_1),
    .O_14_2_2(n97_O_14_2_2),
    .O_15_0_0(n97_O_15_0_0),
    .O_15_0_1(n97_O_15_0_1),
    .O_15_0_2(n97_O_15_0_2),
    .O_15_1_0(n97_O_15_1_0),
    .O_15_1_1(n97_O_15_1_1),
    .O_15_1_2(n97_O_15_1_2),
    .O_15_2_0(n97_O_15_2_0),
    .O_15_2_1(n97_O_15_2_1),
    .O_15_2_2(n97_O_15_2_2)
  );
  MapT_6 n106 ( // @[Top.scala 147:22]
    .valid_up(n106_valid_up),
    .valid_down(n106_valid_down),
    .I_0_0_0(n106_I_0_0_0),
    .I_0_0_1(n106_I_0_0_1),
    .I_0_0_2(n106_I_0_0_2),
    .I_0_1_0(n106_I_0_1_0),
    .I_0_1_1(n106_I_0_1_1),
    .I_0_1_2(n106_I_0_1_2),
    .I_0_2_0(n106_I_0_2_0),
    .I_0_2_1(n106_I_0_2_1),
    .I_0_2_2(n106_I_0_2_2),
    .I_1_0_0(n106_I_1_0_0),
    .I_1_0_1(n106_I_1_0_1),
    .I_1_0_2(n106_I_1_0_2),
    .I_1_1_0(n106_I_1_1_0),
    .I_1_1_1(n106_I_1_1_1),
    .I_1_1_2(n106_I_1_1_2),
    .I_1_2_0(n106_I_1_2_0),
    .I_1_2_1(n106_I_1_2_1),
    .I_1_2_2(n106_I_1_2_2),
    .I_2_0_0(n106_I_2_0_0),
    .I_2_0_1(n106_I_2_0_1),
    .I_2_0_2(n106_I_2_0_2),
    .I_2_1_0(n106_I_2_1_0),
    .I_2_1_1(n106_I_2_1_1),
    .I_2_1_2(n106_I_2_1_2),
    .I_2_2_0(n106_I_2_2_0),
    .I_2_2_1(n106_I_2_2_1),
    .I_2_2_2(n106_I_2_2_2),
    .I_3_0_0(n106_I_3_0_0),
    .I_3_0_1(n106_I_3_0_1),
    .I_3_0_2(n106_I_3_0_2),
    .I_3_1_0(n106_I_3_1_0),
    .I_3_1_1(n106_I_3_1_1),
    .I_3_1_2(n106_I_3_1_2),
    .I_3_2_0(n106_I_3_2_0),
    .I_3_2_1(n106_I_3_2_1),
    .I_3_2_2(n106_I_3_2_2),
    .I_4_0_0(n106_I_4_0_0),
    .I_4_0_1(n106_I_4_0_1),
    .I_4_0_2(n106_I_4_0_2),
    .I_4_1_0(n106_I_4_1_0),
    .I_4_1_1(n106_I_4_1_1),
    .I_4_1_2(n106_I_4_1_2),
    .I_4_2_0(n106_I_4_2_0),
    .I_4_2_1(n106_I_4_2_1),
    .I_4_2_2(n106_I_4_2_2),
    .I_5_0_0(n106_I_5_0_0),
    .I_5_0_1(n106_I_5_0_1),
    .I_5_0_2(n106_I_5_0_2),
    .I_5_1_0(n106_I_5_1_0),
    .I_5_1_1(n106_I_5_1_1),
    .I_5_1_2(n106_I_5_1_2),
    .I_5_2_0(n106_I_5_2_0),
    .I_5_2_1(n106_I_5_2_1),
    .I_5_2_2(n106_I_5_2_2),
    .I_6_0_0(n106_I_6_0_0),
    .I_6_0_1(n106_I_6_0_1),
    .I_6_0_2(n106_I_6_0_2),
    .I_6_1_0(n106_I_6_1_0),
    .I_6_1_1(n106_I_6_1_1),
    .I_6_1_2(n106_I_6_1_2),
    .I_6_2_0(n106_I_6_2_0),
    .I_6_2_1(n106_I_6_2_1),
    .I_6_2_2(n106_I_6_2_2),
    .I_7_0_0(n106_I_7_0_0),
    .I_7_0_1(n106_I_7_0_1),
    .I_7_0_2(n106_I_7_0_2),
    .I_7_1_0(n106_I_7_1_0),
    .I_7_1_1(n106_I_7_1_1),
    .I_7_1_2(n106_I_7_1_2),
    .I_7_2_0(n106_I_7_2_0),
    .I_7_2_1(n106_I_7_2_1),
    .I_7_2_2(n106_I_7_2_2),
    .I_8_0_0(n106_I_8_0_0),
    .I_8_0_1(n106_I_8_0_1),
    .I_8_0_2(n106_I_8_0_2),
    .I_8_1_0(n106_I_8_1_0),
    .I_8_1_1(n106_I_8_1_1),
    .I_8_1_2(n106_I_8_1_2),
    .I_8_2_0(n106_I_8_2_0),
    .I_8_2_1(n106_I_8_2_1),
    .I_8_2_2(n106_I_8_2_2),
    .I_9_0_0(n106_I_9_0_0),
    .I_9_0_1(n106_I_9_0_1),
    .I_9_0_2(n106_I_9_0_2),
    .I_9_1_0(n106_I_9_1_0),
    .I_9_1_1(n106_I_9_1_1),
    .I_9_1_2(n106_I_9_1_2),
    .I_9_2_0(n106_I_9_2_0),
    .I_9_2_1(n106_I_9_2_1),
    .I_9_2_2(n106_I_9_2_2),
    .I_10_0_0(n106_I_10_0_0),
    .I_10_0_1(n106_I_10_0_1),
    .I_10_0_2(n106_I_10_0_2),
    .I_10_1_0(n106_I_10_1_0),
    .I_10_1_1(n106_I_10_1_1),
    .I_10_1_2(n106_I_10_1_2),
    .I_10_2_0(n106_I_10_2_0),
    .I_10_2_1(n106_I_10_2_1),
    .I_10_2_2(n106_I_10_2_2),
    .I_11_0_0(n106_I_11_0_0),
    .I_11_0_1(n106_I_11_0_1),
    .I_11_0_2(n106_I_11_0_2),
    .I_11_1_0(n106_I_11_1_0),
    .I_11_1_1(n106_I_11_1_1),
    .I_11_1_2(n106_I_11_1_2),
    .I_11_2_0(n106_I_11_2_0),
    .I_11_2_1(n106_I_11_2_1),
    .I_11_2_2(n106_I_11_2_2),
    .I_12_0_0(n106_I_12_0_0),
    .I_12_0_1(n106_I_12_0_1),
    .I_12_0_2(n106_I_12_0_2),
    .I_12_1_0(n106_I_12_1_0),
    .I_12_1_1(n106_I_12_1_1),
    .I_12_1_2(n106_I_12_1_2),
    .I_12_2_0(n106_I_12_2_0),
    .I_12_2_1(n106_I_12_2_1),
    .I_12_2_2(n106_I_12_2_2),
    .I_13_0_0(n106_I_13_0_0),
    .I_13_0_1(n106_I_13_0_1),
    .I_13_0_2(n106_I_13_0_2),
    .I_13_1_0(n106_I_13_1_0),
    .I_13_1_1(n106_I_13_1_1),
    .I_13_1_2(n106_I_13_1_2),
    .I_13_2_0(n106_I_13_2_0),
    .I_13_2_1(n106_I_13_2_1),
    .I_13_2_2(n106_I_13_2_2),
    .I_14_0_0(n106_I_14_0_0),
    .I_14_0_1(n106_I_14_0_1),
    .I_14_0_2(n106_I_14_0_2),
    .I_14_1_0(n106_I_14_1_0),
    .I_14_1_1(n106_I_14_1_1),
    .I_14_1_2(n106_I_14_1_2),
    .I_14_2_0(n106_I_14_2_0),
    .I_14_2_1(n106_I_14_2_1),
    .I_14_2_2(n106_I_14_2_2),
    .I_15_0_0(n106_I_15_0_0),
    .I_15_0_1(n106_I_15_0_1),
    .I_15_0_2(n106_I_15_0_2),
    .I_15_1_0(n106_I_15_1_0),
    .I_15_1_1(n106_I_15_1_1),
    .I_15_1_2(n106_I_15_1_2),
    .I_15_2_0(n106_I_15_2_0),
    .I_15_2_1(n106_I_15_2_1),
    .I_15_2_2(n106_I_15_2_2),
    .O_0_0_0_0(n106_O_0_0_0_0),
    .O_0_0_0_1(n106_O_0_0_0_1),
    .O_0_0_0_2(n106_O_0_0_0_2),
    .O_0_0_1_0(n106_O_0_0_1_0),
    .O_0_0_1_1(n106_O_0_0_1_1),
    .O_0_0_1_2(n106_O_0_0_1_2),
    .O_0_0_2_0(n106_O_0_0_2_0),
    .O_0_0_2_1(n106_O_0_0_2_1),
    .O_0_0_2_2(n106_O_0_0_2_2),
    .O_1_0_0_0(n106_O_1_0_0_0),
    .O_1_0_0_1(n106_O_1_0_0_1),
    .O_1_0_0_2(n106_O_1_0_0_2),
    .O_1_0_1_0(n106_O_1_0_1_0),
    .O_1_0_1_1(n106_O_1_0_1_1),
    .O_1_0_1_2(n106_O_1_0_1_2),
    .O_1_0_2_0(n106_O_1_0_2_0),
    .O_1_0_2_1(n106_O_1_0_2_1),
    .O_1_0_2_2(n106_O_1_0_2_2),
    .O_2_0_0_0(n106_O_2_0_0_0),
    .O_2_0_0_1(n106_O_2_0_0_1),
    .O_2_0_0_2(n106_O_2_0_0_2),
    .O_2_0_1_0(n106_O_2_0_1_0),
    .O_2_0_1_1(n106_O_2_0_1_1),
    .O_2_0_1_2(n106_O_2_0_1_2),
    .O_2_0_2_0(n106_O_2_0_2_0),
    .O_2_0_2_1(n106_O_2_0_2_1),
    .O_2_0_2_2(n106_O_2_0_2_2),
    .O_3_0_0_0(n106_O_3_0_0_0),
    .O_3_0_0_1(n106_O_3_0_0_1),
    .O_3_0_0_2(n106_O_3_0_0_2),
    .O_3_0_1_0(n106_O_3_0_1_0),
    .O_3_0_1_1(n106_O_3_0_1_1),
    .O_3_0_1_2(n106_O_3_0_1_2),
    .O_3_0_2_0(n106_O_3_0_2_0),
    .O_3_0_2_1(n106_O_3_0_2_1),
    .O_3_0_2_2(n106_O_3_0_2_2),
    .O_4_0_0_0(n106_O_4_0_0_0),
    .O_4_0_0_1(n106_O_4_0_0_1),
    .O_4_0_0_2(n106_O_4_0_0_2),
    .O_4_0_1_0(n106_O_4_0_1_0),
    .O_4_0_1_1(n106_O_4_0_1_1),
    .O_4_0_1_2(n106_O_4_0_1_2),
    .O_4_0_2_0(n106_O_4_0_2_0),
    .O_4_0_2_1(n106_O_4_0_2_1),
    .O_4_0_2_2(n106_O_4_0_2_2),
    .O_5_0_0_0(n106_O_5_0_0_0),
    .O_5_0_0_1(n106_O_5_0_0_1),
    .O_5_0_0_2(n106_O_5_0_0_2),
    .O_5_0_1_0(n106_O_5_0_1_0),
    .O_5_0_1_1(n106_O_5_0_1_1),
    .O_5_0_1_2(n106_O_5_0_1_2),
    .O_5_0_2_0(n106_O_5_0_2_0),
    .O_5_0_2_1(n106_O_5_0_2_1),
    .O_5_0_2_2(n106_O_5_0_2_2),
    .O_6_0_0_0(n106_O_6_0_0_0),
    .O_6_0_0_1(n106_O_6_0_0_1),
    .O_6_0_0_2(n106_O_6_0_0_2),
    .O_6_0_1_0(n106_O_6_0_1_0),
    .O_6_0_1_1(n106_O_6_0_1_1),
    .O_6_0_1_2(n106_O_6_0_1_2),
    .O_6_0_2_0(n106_O_6_0_2_0),
    .O_6_0_2_1(n106_O_6_0_2_1),
    .O_6_0_2_2(n106_O_6_0_2_2),
    .O_7_0_0_0(n106_O_7_0_0_0),
    .O_7_0_0_1(n106_O_7_0_0_1),
    .O_7_0_0_2(n106_O_7_0_0_2),
    .O_7_0_1_0(n106_O_7_0_1_0),
    .O_7_0_1_1(n106_O_7_0_1_1),
    .O_7_0_1_2(n106_O_7_0_1_2),
    .O_7_0_2_0(n106_O_7_0_2_0),
    .O_7_0_2_1(n106_O_7_0_2_1),
    .O_7_0_2_2(n106_O_7_0_2_2),
    .O_8_0_0_0(n106_O_8_0_0_0),
    .O_8_0_0_1(n106_O_8_0_0_1),
    .O_8_0_0_2(n106_O_8_0_0_2),
    .O_8_0_1_0(n106_O_8_0_1_0),
    .O_8_0_1_1(n106_O_8_0_1_1),
    .O_8_0_1_2(n106_O_8_0_1_2),
    .O_8_0_2_0(n106_O_8_0_2_0),
    .O_8_0_2_1(n106_O_8_0_2_1),
    .O_8_0_2_2(n106_O_8_0_2_2),
    .O_9_0_0_0(n106_O_9_0_0_0),
    .O_9_0_0_1(n106_O_9_0_0_1),
    .O_9_0_0_2(n106_O_9_0_0_2),
    .O_9_0_1_0(n106_O_9_0_1_0),
    .O_9_0_1_1(n106_O_9_0_1_1),
    .O_9_0_1_2(n106_O_9_0_1_2),
    .O_9_0_2_0(n106_O_9_0_2_0),
    .O_9_0_2_1(n106_O_9_0_2_1),
    .O_9_0_2_2(n106_O_9_0_2_2),
    .O_10_0_0_0(n106_O_10_0_0_0),
    .O_10_0_0_1(n106_O_10_0_0_1),
    .O_10_0_0_2(n106_O_10_0_0_2),
    .O_10_0_1_0(n106_O_10_0_1_0),
    .O_10_0_1_1(n106_O_10_0_1_1),
    .O_10_0_1_2(n106_O_10_0_1_2),
    .O_10_0_2_0(n106_O_10_0_2_0),
    .O_10_0_2_1(n106_O_10_0_2_1),
    .O_10_0_2_2(n106_O_10_0_2_2),
    .O_11_0_0_0(n106_O_11_0_0_0),
    .O_11_0_0_1(n106_O_11_0_0_1),
    .O_11_0_0_2(n106_O_11_0_0_2),
    .O_11_0_1_0(n106_O_11_0_1_0),
    .O_11_0_1_1(n106_O_11_0_1_1),
    .O_11_0_1_2(n106_O_11_0_1_2),
    .O_11_0_2_0(n106_O_11_0_2_0),
    .O_11_0_2_1(n106_O_11_0_2_1),
    .O_11_0_2_2(n106_O_11_0_2_2),
    .O_12_0_0_0(n106_O_12_0_0_0),
    .O_12_0_0_1(n106_O_12_0_0_1),
    .O_12_0_0_2(n106_O_12_0_0_2),
    .O_12_0_1_0(n106_O_12_0_1_0),
    .O_12_0_1_1(n106_O_12_0_1_1),
    .O_12_0_1_2(n106_O_12_0_1_2),
    .O_12_0_2_0(n106_O_12_0_2_0),
    .O_12_0_2_1(n106_O_12_0_2_1),
    .O_12_0_2_2(n106_O_12_0_2_2),
    .O_13_0_0_0(n106_O_13_0_0_0),
    .O_13_0_0_1(n106_O_13_0_0_1),
    .O_13_0_0_2(n106_O_13_0_0_2),
    .O_13_0_1_0(n106_O_13_0_1_0),
    .O_13_0_1_1(n106_O_13_0_1_1),
    .O_13_0_1_2(n106_O_13_0_1_2),
    .O_13_0_2_0(n106_O_13_0_2_0),
    .O_13_0_2_1(n106_O_13_0_2_1),
    .O_13_0_2_2(n106_O_13_0_2_2),
    .O_14_0_0_0(n106_O_14_0_0_0),
    .O_14_0_0_1(n106_O_14_0_0_1),
    .O_14_0_0_2(n106_O_14_0_0_2),
    .O_14_0_1_0(n106_O_14_0_1_0),
    .O_14_0_1_1(n106_O_14_0_1_1),
    .O_14_0_1_2(n106_O_14_0_1_2),
    .O_14_0_2_0(n106_O_14_0_2_0),
    .O_14_0_2_1(n106_O_14_0_2_1),
    .O_14_0_2_2(n106_O_14_0_2_2),
    .O_15_0_0_0(n106_O_15_0_0_0),
    .O_15_0_0_1(n106_O_15_0_0_1),
    .O_15_0_0_2(n106_O_15_0_0_2),
    .O_15_0_1_0(n106_O_15_0_1_0),
    .O_15_0_1_1(n106_O_15_0_1_1),
    .O_15_0_1_2(n106_O_15_0_1_2),
    .O_15_0_2_0(n106_O_15_0_2_0),
    .O_15_0_2_1(n106_O_15_0_2_1),
    .O_15_0_2_2(n106_O_15_0_2_2)
  );
  MapT_7 n113 ( // @[Top.scala 150:22]
    .valid_up(n113_valid_up),
    .valid_down(n113_valid_down),
    .I_0_0_0_0(n113_I_0_0_0_0),
    .I_0_0_0_1(n113_I_0_0_0_1),
    .I_0_0_0_2(n113_I_0_0_0_2),
    .I_0_0_1_0(n113_I_0_0_1_0),
    .I_0_0_1_1(n113_I_0_0_1_1),
    .I_0_0_1_2(n113_I_0_0_1_2),
    .I_0_0_2_0(n113_I_0_0_2_0),
    .I_0_0_2_1(n113_I_0_0_2_1),
    .I_0_0_2_2(n113_I_0_0_2_2),
    .I_1_0_0_0(n113_I_1_0_0_0),
    .I_1_0_0_1(n113_I_1_0_0_1),
    .I_1_0_0_2(n113_I_1_0_0_2),
    .I_1_0_1_0(n113_I_1_0_1_0),
    .I_1_0_1_1(n113_I_1_0_1_1),
    .I_1_0_1_2(n113_I_1_0_1_2),
    .I_1_0_2_0(n113_I_1_0_2_0),
    .I_1_0_2_1(n113_I_1_0_2_1),
    .I_1_0_2_2(n113_I_1_0_2_2),
    .I_2_0_0_0(n113_I_2_0_0_0),
    .I_2_0_0_1(n113_I_2_0_0_1),
    .I_2_0_0_2(n113_I_2_0_0_2),
    .I_2_0_1_0(n113_I_2_0_1_0),
    .I_2_0_1_1(n113_I_2_0_1_1),
    .I_2_0_1_2(n113_I_2_0_1_2),
    .I_2_0_2_0(n113_I_2_0_2_0),
    .I_2_0_2_1(n113_I_2_0_2_1),
    .I_2_0_2_2(n113_I_2_0_2_2),
    .I_3_0_0_0(n113_I_3_0_0_0),
    .I_3_0_0_1(n113_I_3_0_0_1),
    .I_3_0_0_2(n113_I_3_0_0_2),
    .I_3_0_1_0(n113_I_3_0_1_0),
    .I_3_0_1_1(n113_I_3_0_1_1),
    .I_3_0_1_2(n113_I_3_0_1_2),
    .I_3_0_2_0(n113_I_3_0_2_0),
    .I_3_0_2_1(n113_I_3_0_2_1),
    .I_3_0_2_2(n113_I_3_0_2_2),
    .I_4_0_0_0(n113_I_4_0_0_0),
    .I_4_0_0_1(n113_I_4_0_0_1),
    .I_4_0_0_2(n113_I_4_0_0_2),
    .I_4_0_1_0(n113_I_4_0_1_0),
    .I_4_0_1_1(n113_I_4_0_1_1),
    .I_4_0_1_2(n113_I_4_0_1_2),
    .I_4_0_2_0(n113_I_4_0_2_0),
    .I_4_0_2_1(n113_I_4_0_2_1),
    .I_4_0_2_2(n113_I_4_0_2_2),
    .I_5_0_0_0(n113_I_5_0_0_0),
    .I_5_0_0_1(n113_I_5_0_0_1),
    .I_5_0_0_2(n113_I_5_0_0_2),
    .I_5_0_1_0(n113_I_5_0_1_0),
    .I_5_0_1_1(n113_I_5_0_1_1),
    .I_5_0_1_2(n113_I_5_0_1_2),
    .I_5_0_2_0(n113_I_5_0_2_0),
    .I_5_0_2_1(n113_I_5_0_2_1),
    .I_5_0_2_2(n113_I_5_0_2_2),
    .I_6_0_0_0(n113_I_6_0_0_0),
    .I_6_0_0_1(n113_I_6_0_0_1),
    .I_6_0_0_2(n113_I_6_0_0_2),
    .I_6_0_1_0(n113_I_6_0_1_0),
    .I_6_0_1_1(n113_I_6_0_1_1),
    .I_6_0_1_2(n113_I_6_0_1_2),
    .I_6_0_2_0(n113_I_6_0_2_0),
    .I_6_0_2_1(n113_I_6_0_2_1),
    .I_6_0_2_2(n113_I_6_0_2_2),
    .I_7_0_0_0(n113_I_7_0_0_0),
    .I_7_0_0_1(n113_I_7_0_0_1),
    .I_7_0_0_2(n113_I_7_0_0_2),
    .I_7_0_1_0(n113_I_7_0_1_0),
    .I_7_0_1_1(n113_I_7_0_1_1),
    .I_7_0_1_2(n113_I_7_0_1_2),
    .I_7_0_2_0(n113_I_7_0_2_0),
    .I_7_0_2_1(n113_I_7_0_2_1),
    .I_7_0_2_2(n113_I_7_0_2_2),
    .I_8_0_0_0(n113_I_8_0_0_0),
    .I_8_0_0_1(n113_I_8_0_0_1),
    .I_8_0_0_2(n113_I_8_0_0_2),
    .I_8_0_1_0(n113_I_8_0_1_0),
    .I_8_0_1_1(n113_I_8_0_1_1),
    .I_8_0_1_2(n113_I_8_0_1_2),
    .I_8_0_2_0(n113_I_8_0_2_0),
    .I_8_0_2_1(n113_I_8_0_2_1),
    .I_8_0_2_2(n113_I_8_0_2_2),
    .I_9_0_0_0(n113_I_9_0_0_0),
    .I_9_0_0_1(n113_I_9_0_0_1),
    .I_9_0_0_2(n113_I_9_0_0_2),
    .I_9_0_1_0(n113_I_9_0_1_0),
    .I_9_0_1_1(n113_I_9_0_1_1),
    .I_9_0_1_2(n113_I_9_0_1_2),
    .I_9_0_2_0(n113_I_9_0_2_0),
    .I_9_0_2_1(n113_I_9_0_2_1),
    .I_9_0_2_2(n113_I_9_0_2_2),
    .I_10_0_0_0(n113_I_10_0_0_0),
    .I_10_0_0_1(n113_I_10_0_0_1),
    .I_10_0_0_2(n113_I_10_0_0_2),
    .I_10_0_1_0(n113_I_10_0_1_0),
    .I_10_0_1_1(n113_I_10_0_1_1),
    .I_10_0_1_2(n113_I_10_0_1_2),
    .I_10_0_2_0(n113_I_10_0_2_0),
    .I_10_0_2_1(n113_I_10_0_2_1),
    .I_10_0_2_2(n113_I_10_0_2_2),
    .I_11_0_0_0(n113_I_11_0_0_0),
    .I_11_0_0_1(n113_I_11_0_0_1),
    .I_11_0_0_2(n113_I_11_0_0_2),
    .I_11_0_1_0(n113_I_11_0_1_0),
    .I_11_0_1_1(n113_I_11_0_1_1),
    .I_11_0_1_2(n113_I_11_0_1_2),
    .I_11_0_2_0(n113_I_11_0_2_0),
    .I_11_0_2_1(n113_I_11_0_2_1),
    .I_11_0_2_2(n113_I_11_0_2_2),
    .I_12_0_0_0(n113_I_12_0_0_0),
    .I_12_0_0_1(n113_I_12_0_0_1),
    .I_12_0_0_2(n113_I_12_0_0_2),
    .I_12_0_1_0(n113_I_12_0_1_0),
    .I_12_0_1_1(n113_I_12_0_1_1),
    .I_12_0_1_2(n113_I_12_0_1_2),
    .I_12_0_2_0(n113_I_12_0_2_0),
    .I_12_0_2_1(n113_I_12_0_2_1),
    .I_12_0_2_2(n113_I_12_0_2_2),
    .I_13_0_0_0(n113_I_13_0_0_0),
    .I_13_0_0_1(n113_I_13_0_0_1),
    .I_13_0_0_2(n113_I_13_0_0_2),
    .I_13_0_1_0(n113_I_13_0_1_0),
    .I_13_0_1_1(n113_I_13_0_1_1),
    .I_13_0_1_2(n113_I_13_0_1_2),
    .I_13_0_2_0(n113_I_13_0_2_0),
    .I_13_0_2_1(n113_I_13_0_2_1),
    .I_13_0_2_2(n113_I_13_0_2_2),
    .I_14_0_0_0(n113_I_14_0_0_0),
    .I_14_0_0_1(n113_I_14_0_0_1),
    .I_14_0_0_2(n113_I_14_0_0_2),
    .I_14_0_1_0(n113_I_14_0_1_0),
    .I_14_0_1_1(n113_I_14_0_1_1),
    .I_14_0_1_2(n113_I_14_0_1_2),
    .I_14_0_2_0(n113_I_14_0_2_0),
    .I_14_0_2_1(n113_I_14_0_2_1),
    .I_14_0_2_2(n113_I_14_0_2_2),
    .I_15_0_0_0(n113_I_15_0_0_0),
    .I_15_0_0_1(n113_I_15_0_0_1),
    .I_15_0_0_2(n113_I_15_0_0_2),
    .I_15_0_1_0(n113_I_15_0_1_0),
    .I_15_0_1_1(n113_I_15_0_1_1),
    .I_15_0_1_2(n113_I_15_0_1_2),
    .I_15_0_2_0(n113_I_15_0_2_0),
    .I_15_0_2_1(n113_I_15_0_2_1),
    .I_15_0_2_2(n113_I_15_0_2_2),
    .O_0_0_0(n113_O_0_0_0),
    .O_0_0_1(n113_O_0_0_1),
    .O_0_0_2(n113_O_0_0_2),
    .O_0_1_0(n113_O_0_1_0),
    .O_0_1_1(n113_O_0_1_1),
    .O_0_1_2(n113_O_0_1_2),
    .O_0_2_0(n113_O_0_2_0),
    .O_0_2_1(n113_O_0_2_1),
    .O_0_2_2(n113_O_0_2_2),
    .O_1_0_0(n113_O_1_0_0),
    .O_1_0_1(n113_O_1_0_1),
    .O_1_0_2(n113_O_1_0_2),
    .O_1_1_0(n113_O_1_1_0),
    .O_1_1_1(n113_O_1_1_1),
    .O_1_1_2(n113_O_1_1_2),
    .O_1_2_0(n113_O_1_2_0),
    .O_1_2_1(n113_O_1_2_1),
    .O_1_2_2(n113_O_1_2_2),
    .O_2_0_0(n113_O_2_0_0),
    .O_2_0_1(n113_O_2_0_1),
    .O_2_0_2(n113_O_2_0_2),
    .O_2_1_0(n113_O_2_1_0),
    .O_2_1_1(n113_O_2_1_1),
    .O_2_1_2(n113_O_2_1_2),
    .O_2_2_0(n113_O_2_2_0),
    .O_2_2_1(n113_O_2_2_1),
    .O_2_2_2(n113_O_2_2_2),
    .O_3_0_0(n113_O_3_0_0),
    .O_3_0_1(n113_O_3_0_1),
    .O_3_0_2(n113_O_3_0_2),
    .O_3_1_0(n113_O_3_1_0),
    .O_3_1_1(n113_O_3_1_1),
    .O_3_1_2(n113_O_3_1_2),
    .O_3_2_0(n113_O_3_2_0),
    .O_3_2_1(n113_O_3_2_1),
    .O_3_2_2(n113_O_3_2_2),
    .O_4_0_0(n113_O_4_0_0),
    .O_4_0_1(n113_O_4_0_1),
    .O_4_0_2(n113_O_4_0_2),
    .O_4_1_0(n113_O_4_1_0),
    .O_4_1_1(n113_O_4_1_1),
    .O_4_1_2(n113_O_4_1_2),
    .O_4_2_0(n113_O_4_2_0),
    .O_4_2_1(n113_O_4_2_1),
    .O_4_2_2(n113_O_4_2_2),
    .O_5_0_0(n113_O_5_0_0),
    .O_5_0_1(n113_O_5_0_1),
    .O_5_0_2(n113_O_5_0_2),
    .O_5_1_0(n113_O_5_1_0),
    .O_5_1_1(n113_O_5_1_1),
    .O_5_1_2(n113_O_5_1_2),
    .O_5_2_0(n113_O_5_2_0),
    .O_5_2_1(n113_O_5_2_1),
    .O_5_2_2(n113_O_5_2_2),
    .O_6_0_0(n113_O_6_0_0),
    .O_6_0_1(n113_O_6_0_1),
    .O_6_0_2(n113_O_6_0_2),
    .O_6_1_0(n113_O_6_1_0),
    .O_6_1_1(n113_O_6_1_1),
    .O_6_1_2(n113_O_6_1_2),
    .O_6_2_0(n113_O_6_2_0),
    .O_6_2_1(n113_O_6_2_1),
    .O_6_2_2(n113_O_6_2_2),
    .O_7_0_0(n113_O_7_0_0),
    .O_7_0_1(n113_O_7_0_1),
    .O_7_0_2(n113_O_7_0_2),
    .O_7_1_0(n113_O_7_1_0),
    .O_7_1_1(n113_O_7_1_1),
    .O_7_1_2(n113_O_7_1_2),
    .O_7_2_0(n113_O_7_2_0),
    .O_7_2_1(n113_O_7_2_1),
    .O_7_2_2(n113_O_7_2_2),
    .O_8_0_0(n113_O_8_0_0),
    .O_8_0_1(n113_O_8_0_1),
    .O_8_0_2(n113_O_8_0_2),
    .O_8_1_0(n113_O_8_1_0),
    .O_8_1_1(n113_O_8_1_1),
    .O_8_1_2(n113_O_8_1_2),
    .O_8_2_0(n113_O_8_2_0),
    .O_8_2_1(n113_O_8_2_1),
    .O_8_2_2(n113_O_8_2_2),
    .O_9_0_0(n113_O_9_0_0),
    .O_9_0_1(n113_O_9_0_1),
    .O_9_0_2(n113_O_9_0_2),
    .O_9_1_0(n113_O_9_1_0),
    .O_9_1_1(n113_O_9_1_1),
    .O_9_1_2(n113_O_9_1_2),
    .O_9_2_0(n113_O_9_2_0),
    .O_9_2_1(n113_O_9_2_1),
    .O_9_2_2(n113_O_9_2_2),
    .O_10_0_0(n113_O_10_0_0),
    .O_10_0_1(n113_O_10_0_1),
    .O_10_0_2(n113_O_10_0_2),
    .O_10_1_0(n113_O_10_1_0),
    .O_10_1_1(n113_O_10_1_1),
    .O_10_1_2(n113_O_10_1_2),
    .O_10_2_0(n113_O_10_2_0),
    .O_10_2_1(n113_O_10_2_1),
    .O_10_2_2(n113_O_10_2_2),
    .O_11_0_0(n113_O_11_0_0),
    .O_11_0_1(n113_O_11_0_1),
    .O_11_0_2(n113_O_11_0_2),
    .O_11_1_0(n113_O_11_1_0),
    .O_11_1_1(n113_O_11_1_1),
    .O_11_1_2(n113_O_11_1_2),
    .O_11_2_0(n113_O_11_2_0),
    .O_11_2_1(n113_O_11_2_1),
    .O_11_2_2(n113_O_11_2_2),
    .O_12_0_0(n113_O_12_0_0),
    .O_12_0_1(n113_O_12_0_1),
    .O_12_0_2(n113_O_12_0_2),
    .O_12_1_0(n113_O_12_1_0),
    .O_12_1_1(n113_O_12_1_1),
    .O_12_1_2(n113_O_12_1_2),
    .O_12_2_0(n113_O_12_2_0),
    .O_12_2_1(n113_O_12_2_1),
    .O_12_2_2(n113_O_12_2_2),
    .O_13_0_0(n113_O_13_0_0),
    .O_13_0_1(n113_O_13_0_1),
    .O_13_0_2(n113_O_13_0_2),
    .O_13_1_0(n113_O_13_1_0),
    .O_13_1_1(n113_O_13_1_1),
    .O_13_1_2(n113_O_13_1_2),
    .O_13_2_0(n113_O_13_2_0),
    .O_13_2_1(n113_O_13_2_1),
    .O_13_2_2(n113_O_13_2_2),
    .O_14_0_0(n113_O_14_0_0),
    .O_14_0_1(n113_O_14_0_1),
    .O_14_0_2(n113_O_14_0_2),
    .O_14_1_0(n113_O_14_1_0),
    .O_14_1_1(n113_O_14_1_1),
    .O_14_1_2(n113_O_14_1_2),
    .O_14_2_0(n113_O_14_2_0),
    .O_14_2_1(n113_O_14_2_1),
    .O_14_2_2(n113_O_14_2_2),
    .O_15_0_0(n113_O_15_0_0),
    .O_15_0_1(n113_O_15_0_1),
    .O_15_0_2(n113_O_15_0_2),
    .O_15_1_0(n113_O_15_1_0),
    .O_15_1_1(n113_O_15_1_1),
    .O_15_1_2(n113_O_15_1_2),
    .O_15_2_0(n113_O_15_2_0),
    .O_15_2_1(n113_O_15_2_1),
    .O_15_2_2(n113_O_15_2_2)
  );
  MapT_8 n155 ( // @[Top.scala 153:22]
    .clock(n155_clock),
    .reset(n155_reset),
    .valid_up(n155_valid_up),
    .valid_down(n155_valid_down),
    .I_0_0_0(n155_I_0_0_0),
    .I_0_0_1(n155_I_0_0_1),
    .I_0_0_2(n155_I_0_0_2),
    .I_0_1_0(n155_I_0_1_0),
    .I_0_1_1(n155_I_0_1_1),
    .I_0_1_2(n155_I_0_1_2),
    .I_0_2_0(n155_I_0_2_0),
    .I_0_2_1(n155_I_0_2_1),
    .I_0_2_2(n155_I_0_2_2),
    .I_1_0_0(n155_I_1_0_0),
    .I_1_0_1(n155_I_1_0_1),
    .I_1_0_2(n155_I_1_0_2),
    .I_1_1_0(n155_I_1_1_0),
    .I_1_1_1(n155_I_1_1_1),
    .I_1_1_2(n155_I_1_1_2),
    .I_1_2_0(n155_I_1_2_0),
    .I_1_2_1(n155_I_1_2_1),
    .I_1_2_2(n155_I_1_2_2),
    .I_2_0_0(n155_I_2_0_0),
    .I_2_0_1(n155_I_2_0_1),
    .I_2_0_2(n155_I_2_0_2),
    .I_2_1_0(n155_I_2_1_0),
    .I_2_1_1(n155_I_2_1_1),
    .I_2_1_2(n155_I_2_1_2),
    .I_2_2_0(n155_I_2_2_0),
    .I_2_2_1(n155_I_2_2_1),
    .I_2_2_2(n155_I_2_2_2),
    .I_3_0_0(n155_I_3_0_0),
    .I_3_0_1(n155_I_3_0_1),
    .I_3_0_2(n155_I_3_0_2),
    .I_3_1_0(n155_I_3_1_0),
    .I_3_1_1(n155_I_3_1_1),
    .I_3_1_2(n155_I_3_1_2),
    .I_3_2_0(n155_I_3_2_0),
    .I_3_2_1(n155_I_3_2_1),
    .I_3_2_2(n155_I_3_2_2),
    .I_4_0_0(n155_I_4_0_0),
    .I_4_0_1(n155_I_4_0_1),
    .I_4_0_2(n155_I_4_0_2),
    .I_4_1_0(n155_I_4_1_0),
    .I_4_1_1(n155_I_4_1_1),
    .I_4_1_2(n155_I_4_1_2),
    .I_4_2_0(n155_I_4_2_0),
    .I_4_2_1(n155_I_4_2_1),
    .I_4_2_2(n155_I_4_2_2),
    .I_5_0_0(n155_I_5_0_0),
    .I_5_0_1(n155_I_5_0_1),
    .I_5_0_2(n155_I_5_0_2),
    .I_5_1_0(n155_I_5_1_0),
    .I_5_1_1(n155_I_5_1_1),
    .I_5_1_2(n155_I_5_1_2),
    .I_5_2_0(n155_I_5_2_0),
    .I_5_2_1(n155_I_5_2_1),
    .I_5_2_2(n155_I_5_2_2),
    .I_6_0_0(n155_I_6_0_0),
    .I_6_0_1(n155_I_6_0_1),
    .I_6_0_2(n155_I_6_0_2),
    .I_6_1_0(n155_I_6_1_0),
    .I_6_1_1(n155_I_6_1_1),
    .I_6_1_2(n155_I_6_1_2),
    .I_6_2_0(n155_I_6_2_0),
    .I_6_2_1(n155_I_6_2_1),
    .I_6_2_2(n155_I_6_2_2),
    .I_7_0_0(n155_I_7_0_0),
    .I_7_0_1(n155_I_7_0_1),
    .I_7_0_2(n155_I_7_0_2),
    .I_7_1_0(n155_I_7_1_0),
    .I_7_1_1(n155_I_7_1_1),
    .I_7_1_2(n155_I_7_1_2),
    .I_7_2_0(n155_I_7_2_0),
    .I_7_2_1(n155_I_7_2_1),
    .I_7_2_2(n155_I_7_2_2),
    .I_8_0_0(n155_I_8_0_0),
    .I_8_0_1(n155_I_8_0_1),
    .I_8_0_2(n155_I_8_0_2),
    .I_8_1_0(n155_I_8_1_0),
    .I_8_1_1(n155_I_8_1_1),
    .I_8_1_2(n155_I_8_1_2),
    .I_8_2_0(n155_I_8_2_0),
    .I_8_2_1(n155_I_8_2_1),
    .I_8_2_2(n155_I_8_2_2),
    .I_9_0_0(n155_I_9_0_0),
    .I_9_0_1(n155_I_9_0_1),
    .I_9_0_2(n155_I_9_0_2),
    .I_9_1_0(n155_I_9_1_0),
    .I_9_1_1(n155_I_9_1_1),
    .I_9_1_2(n155_I_9_1_2),
    .I_9_2_0(n155_I_9_2_0),
    .I_9_2_1(n155_I_9_2_1),
    .I_9_2_2(n155_I_9_2_2),
    .I_10_0_0(n155_I_10_0_0),
    .I_10_0_1(n155_I_10_0_1),
    .I_10_0_2(n155_I_10_0_2),
    .I_10_1_0(n155_I_10_1_0),
    .I_10_1_1(n155_I_10_1_1),
    .I_10_1_2(n155_I_10_1_2),
    .I_10_2_0(n155_I_10_2_0),
    .I_10_2_1(n155_I_10_2_1),
    .I_10_2_2(n155_I_10_2_2),
    .I_11_0_0(n155_I_11_0_0),
    .I_11_0_1(n155_I_11_0_1),
    .I_11_0_2(n155_I_11_0_2),
    .I_11_1_0(n155_I_11_1_0),
    .I_11_1_1(n155_I_11_1_1),
    .I_11_1_2(n155_I_11_1_2),
    .I_11_2_0(n155_I_11_2_0),
    .I_11_2_1(n155_I_11_2_1),
    .I_11_2_2(n155_I_11_2_2),
    .I_12_0_0(n155_I_12_0_0),
    .I_12_0_1(n155_I_12_0_1),
    .I_12_0_2(n155_I_12_0_2),
    .I_12_1_0(n155_I_12_1_0),
    .I_12_1_1(n155_I_12_1_1),
    .I_12_1_2(n155_I_12_1_2),
    .I_12_2_0(n155_I_12_2_0),
    .I_12_2_1(n155_I_12_2_1),
    .I_12_2_2(n155_I_12_2_2),
    .I_13_0_0(n155_I_13_0_0),
    .I_13_0_1(n155_I_13_0_1),
    .I_13_0_2(n155_I_13_0_2),
    .I_13_1_0(n155_I_13_1_0),
    .I_13_1_1(n155_I_13_1_1),
    .I_13_1_2(n155_I_13_1_2),
    .I_13_2_0(n155_I_13_2_0),
    .I_13_2_1(n155_I_13_2_1),
    .I_13_2_2(n155_I_13_2_2),
    .I_14_0_0(n155_I_14_0_0),
    .I_14_0_1(n155_I_14_0_1),
    .I_14_0_2(n155_I_14_0_2),
    .I_14_1_0(n155_I_14_1_0),
    .I_14_1_1(n155_I_14_1_1),
    .I_14_1_2(n155_I_14_1_2),
    .I_14_2_0(n155_I_14_2_0),
    .I_14_2_1(n155_I_14_2_1),
    .I_14_2_2(n155_I_14_2_2),
    .I_15_0_0(n155_I_15_0_0),
    .I_15_0_1(n155_I_15_0_1),
    .I_15_0_2(n155_I_15_0_2),
    .I_15_1_0(n155_I_15_1_0),
    .I_15_1_1(n155_I_15_1_1),
    .I_15_1_2(n155_I_15_1_2),
    .I_15_2_0(n155_I_15_2_0),
    .I_15_2_1(n155_I_15_2_1),
    .I_15_2_2(n155_I_15_2_2),
    .O_0_0_0(n155_O_0_0_0),
    .O_1_0_0(n155_O_1_0_0),
    .O_2_0_0(n155_O_2_0_0),
    .O_3_0_0(n155_O_3_0_0),
    .O_4_0_0(n155_O_4_0_0),
    .O_5_0_0(n155_O_5_0_0),
    .O_6_0_0(n155_O_6_0_0),
    .O_7_0_0(n155_O_7_0_0),
    .O_8_0_0(n155_O_8_0_0),
    .O_9_0_0(n155_O_9_0_0),
    .O_10_0_0(n155_O_10_0_0),
    .O_11_0_0(n155_O_11_0_0),
    .O_12_0_0(n155_O_12_0_0),
    .O_13_0_0(n155_O_13_0_0),
    .O_14_0_0(n155_O_14_0_0),
    .O_15_0_0(n155_O_15_0_0)
  );
  Passthrough n156 ( // @[Top.scala 156:22]
    .valid_up(n156_valid_up),
    .valid_down(n156_valid_down),
    .I_0_0_0(n156_I_0_0_0),
    .I_1_0_0(n156_I_1_0_0),
    .I_2_0_0(n156_I_2_0_0),
    .I_3_0_0(n156_I_3_0_0),
    .I_4_0_0(n156_I_4_0_0),
    .I_5_0_0(n156_I_5_0_0),
    .I_6_0_0(n156_I_6_0_0),
    .I_7_0_0(n156_I_7_0_0),
    .I_8_0_0(n156_I_8_0_0),
    .I_9_0_0(n156_I_9_0_0),
    .I_10_0_0(n156_I_10_0_0),
    .I_11_0_0(n156_I_11_0_0),
    .I_12_0_0(n156_I_12_0_0),
    .I_13_0_0(n156_I_13_0_0),
    .I_14_0_0(n156_I_14_0_0),
    .I_15_0_0(n156_I_15_0_0),
    .O_0_0(n156_O_0_0),
    .O_1_0(n156_O_1_0),
    .O_2_0(n156_O_2_0),
    .O_3_0(n156_O_3_0),
    .O_4_0(n156_O_4_0),
    .O_5_0(n156_O_5_0),
    .O_6_0(n156_O_6_0),
    .O_7_0(n156_O_7_0),
    .O_8_0(n156_O_8_0),
    .O_9_0(n156_O_9_0),
    .O_10_0(n156_O_10_0),
    .O_11_0(n156_O_11_0),
    .O_12_0(n156_O_12_0),
    .O_13_0(n156_O_13_0),
    .O_14_0(n156_O_14_0),
    .O_15_0(n156_O_15_0)
  );
  Passthrough_1 n157 ( // @[Top.scala 159:22]
    .valid_up(n157_valid_up),
    .valid_down(n157_valid_down),
    .I_0_0(n157_I_0_0),
    .I_1_0(n157_I_1_0),
    .I_2_0(n157_I_2_0),
    .I_3_0(n157_I_3_0),
    .I_4_0(n157_I_4_0),
    .I_5_0(n157_I_5_0),
    .I_6_0(n157_I_6_0),
    .I_7_0(n157_I_7_0),
    .I_8_0(n157_I_8_0),
    .I_9_0(n157_I_9_0),
    .I_10_0(n157_I_10_0),
    .I_11_0(n157_I_11_0),
    .I_12_0(n157_I_12_0),
    .I_13_0(n157_I_13_0),
    .I_14_0(n157_I_14_0),
    .I_15_0(n157_I_15_0),
    .O_0(n157_O_0),
    .O_1(n157_O_1),
    .O_2(n157_O_2),
    .O_3(n157_O_3),
    .O_4(n157_O_4),
    .O_5(n157_O_5),
    .O_6(n157_O_6),
    .O_7(n157_O_7),
    .O_8(n157_O_8),
    .O_9(n157_O_9),
    .O_10(n157_O_10),
    .O_11(n157_O_11),
    .O_12(n157_O_12),
    .O_13(n157_O_13),
    .O_14(n157_O_14),
    .O_15(n157_O_15)
  );
  FIFO n158 ( // @[Top.scala 162:22]
    .clock(n158_clock),
    .reset(n158_reset),
    .valid_up(n158_valid_up),
    .valid_down(n158_valid_down),
    .I_0(n158_I_0),
    .I_1(n158_I_1),
    .I_2(n158_I_2),
    .I_3(n158_I_3),
    .I_4(n158_I_4),
    .I_5(n158_I_5),
    .I_6(n158_I_6),
    .I_7(n158_I_7),
    .I_8(n158_I_8),
    .I_9(n158_I_9),
    .I_10(n158_I_10),
    .I_11(n158_I_11),
    .I_12(n158_I_12),
    .I_13(n158_I_13),
    .I_14(n158_I_14),
    .I_15(n158_I_15),
    .O_0(n158_O_0),
    .O_1(n158_O_1),
    .O_2(n158_O_2),
    .O_3(n158_O_3),
    .O_4(n158_O_4),
    .O_5(n158_O_5),
    .O_6(n158_O_6),
    .O_7(n158_O_7),
    .O_8(n158_O_8),
    .O_9(n158_O_9),
    .O_10(n158_O_10),
    .O_11(n158_O_11),
    .O_12(n158_O_12),
    .O_13(n158_O_13),
    .O_14(n158_O_14),
    .O_15(n158_O_15)
  );
  FIFO n159 ( // @[Top.scala 165:22]
    .clock(n159_clock),
    .reset(n159_reset),
    .valid_up(n159_valid_up),
    .valid_down(n159_valid_down),
    .I_0(n159_I_0),
    .I_1(n159_I_1),
    .I_2(n159_I_2),
    .I_3(n159_I_3),
    .I_4(n159_I_4),
    .I_5(n159_I_5),
    .I_6(n159_I_6),
    .I_7(n159_I_7),
    .I_8(n159_I_8),
    .I_9(n159_I_9),
    .I_10(n159_I_10),
    .I_11(n159_I_11),
    .I_12(n159_I_12),
    .I_13(n159_I_13),
    .I_14(n159_I_14),
    .I_15(n159_I_15),
    .O_0(n159_O_0),
    .O_1(n159_O_1),
    .O_2(n159_O_2),
    .O_3(n159_O_3),
    .O_4(n159_O_4),
    .O_5(n159_O_5),
    .O_6(n159_O_6),
    .O_7(n159_O_7),
    .O_8(n159_O_8),
    .O_9(n159_O_9),
    .O_10(n159_O_10),
    .O_11(n159_O_11),
    .O_12(n159_O_12),
    .O_13(n159_O_13),
    .O_14(n159_O_14),
    .O_15(n159_O_15)
  );
  FIFO n160 ( // @[Top.scala 168:22]
    .clock(n160_clock),
    .reset(n160_reset),
    .valid_up(n160_valid_up),
    .valid_down(n160_valid_down),
    .I_0(n160_I_0),
    .I_1(n160_I_1),
    .I_2(n160_I_2),
    .I_3(n160_I_3),
    .I_4(n160_I_4),
    .I_5(n160_I_5),
    .I_6(n160_I_6),
    .I_7(n160_I_7),
    .I_8(n160_I_8),
    .I_9(n160_I_9),
    .I_10(n160_I_10),
    .I_11(n160_I_11),
    .I_12(n160_I_12),
    .I_13(n160_I_13),
    .I_14(n160_I_14),
    .I_15(n160_I_15),
    .O_0(n160_O_0),
    .O_1(n160_O_1),
    .O_2(n160_O_2),
    .O_3(n160_O_3),
    .O_4(n160_O_4),
    .O_5(n160_O_5),
    .O_6(n160_O_6),
    .O_7(n160_O_7),
    .O_8(n160_O_8),
    .O_9(n160_O_9),
    .O_10(n160_O_10),
    .O_11(n160_O_11),
    .O_12(n160_O_12),
    .O_13(n160_O_13),
    .O_14(n160_O_14),
    .O_15(n160_O_15)
  );
  assign valid_down = n160_valid_down; // @[Top.scala 172:16]
  assign O_0 = n160_O_0; // @[Top.scala 171:7]
  assign O_1 = n160_O_1; // @[Top.scala 171:7]
  assign O_2 = n160_O_2; // @[Top.scala 171:7]
  assign O_3 = n160_O_3; // @[Top.scala 171:7]
  assign O_4 = n160_O_4; // @[Top.scala 171:7]
  assign O_5 = n160_O_5; // @[Top.scala 171:7]
  assign O_6 = n160_O_6; // @[Top.scala 171:7]
  assign O_7 = n160_O_7; // @[Top.scala 171:7]
  assign O_8 = n160_O_8; // @[Top.scala 171:7]
  assign O_9 = n160_O_9; // @[Top.scala 171:7]
  assign O_10 = n160_O_10; // @[Top.scala 171:7]
  assign O_11 = n160_O_11; // @[Top.scala 171:7]
  assign O_12 = n160_O_12; // @[Top.scala 171:7]
  assign O_13 = n160_O_13; // @[Top.scala 171:7]
  assign O_14 = n160_O_14; // @[Top.scala 171:7]
  assign O_15 = n160_O_15; // @[Top.scala 171:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 48:17]
  assign n1_I_0 = I_0; // @[Top.scala 47:10]
  assign n1_I_1 = I_1; // @[Top.scala 47:10]
  assign n1_I_2 = I_2; // @[Top.scala 47:10]
  assign n1_I_3 = I_3; // @[Top.scala 47:10]
  assign n1_I_4 = I_4; // @[Top.scala 47:10]
  assign n1_I_5 = I_5; // @[Top.scala 47:10]
  assign n1_I_6 = I_6; // @[Top.scala 47:10]
  assign n1_I_7 = I_7; // @[Top.scala 47:10]
  assign n1_I_8 = I_8; // @[Top.scala 47:10]
  assign n1_I_9 = I_9; // @[Top.scala 47:10]
  assign n1_I_10 = I_10; // @[Top.scala 47:10]
  assign n1_I_11 = I_11; // @[Top.scala 47:10]
  assign n1_I_12 = I_12; // @[Top.scala 47:10]
  assign n1_I_13 = I_13; // @[Top.scala 47:10]
  assign n1_I_14 = I_14; // @[Top.scala 47:10]
  assign n1_I_15 = I_15; // @[Top.scala 47:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 51:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 50:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 50:10]
  assign n2_I_2 = n1_O_2; // @[Top.scala 50:10]
  assign n2_I_3 = n1_O_3; // @[Top.scala 50:10]
  assign n2_I_4 = n1_O_4; // @[Top.scala 50:10]
  assign n2_I_5 = n1_O_5; // @[Top.scala 50:10]
  assign n2_I_6 = n1_O_6; // @[Top.scala 50:10]
  assign n2_I_7 = n1_O_7; // @[Top.scala 50:10]
  assign n2_I_8 = n1_O_8; // @[Top.scala 50:10]
  assign n2_I_9 = n1_O_9; // @[Top.scala 50:10]
  assign n2_I_10 = n1_O_10; // @[Top.scala 50:10]
  assign n2_I_11 = n1_O_11; // @[Top.scala 50:10]
  assign n2_I_12 = n1_O_12; // @[Top.scala 50:10]
  assign n2_I_13 = n1_O_13; // @[Top.scala 50:10]
  assign n2_I_14 = n1_O_14; // @[Top.scala 50:10]
  assign n2_I_15 = n1_O_15; // @[Top.scala 50:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 54:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 53:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 53:10]
  assign n3_I_2 = n2_O_2; // @[Top.scala 53:10]
  assign n3_I_3 = n2_O_3; // @[Top.scala 53:10]
  assign n3_I_4 = n2_O_4; // @[Top.scala 53:10]
  assign n3_I_5 = n2_O_5; // @[Top.scala 53:10]
  assign n3_I_6 = n2_O_6; // @[Top.scala 53:10]
  assign n3_I_7 = n2_O_7; // @[Top.scala 53:10]
  assign n3_I_8 = n2_O_8; // @[Top.scala 53:10]
  assign n3_I_9 = n2_O_9; // @[Top.scala 53:10]
  assign n3_I_10 = n2_O_10; // @[Top.scala 53:10]
  assign n3_I_11 = n2_O_11; // @[Top.scala 53:10]
  assign n3_I_12 = n2_O_12; // @[Top.scala 53:10]
  assign n3_I_13 = n2_O_13; // @[Top.scala 53:10]
  assign n3_I_14 = n2_O_14; // @[Top.scala 53:10]
  assign n3_I_15 = n2_O_15; // @[Top.scala 53:10]
  assign n4_clock = clock;
  assign n4_reset = reset;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 57:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 56:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 56:10]
  assign n4_I_2 = n3_O_2; // @[Top.scala 56:10]
  assign n4_I_3 = n3_O_3; // @[Top.scala 56:10]
  assign n4_I_4 = n3_O_4; // @[Top.scala 56:10]
  assign n4_I_5 = n3_O_5; // @[Top.scala 56:10]
  assign n4_I_6 = n3_O_6; // @[Top.scala 56:10]
  assign n4_I_7 = n3_O_7; // @[Top.scala 56:10]
  assign n4_I_8 = n3_O_8; // @[Top.scala 56:10]
  assign n4_I_9 = n3_O_9; // @[Top.scala 56:10]
  assign n4_I_10 = n3_O_10; // @[Top.scala 56:10]
  assign n4_I_11 = n3_O_11; // @[Top.scala 56:10]
  assign n4_I_12 = n3_O_12; // @[Top.scala 56:10]
  assign n4_I_13 = n3_O_13; // @[Top.scala 56:10]
  assign n4_I_14 = n3_O_14; // @[Top.scala 56:10]
  assign n4_I_15 = n3_O_15; // @[Top.scala 56:10]
  assign n5_clock = clock;
  assign n5_reset = reset;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 60:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 59:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 59:10]
  assign n5_I_2 = n4_O_2; // @[Top.scala 59:10]
  assign n5_I_3 = n4_O_3; // @[Top.scala 59:10]
  assign n5_I_4 = n4_O_4; // @[Top.scala 59:10]
  assign n5_I_5 = n4_O_5; // @[Top.scala 59:10]
  assign n5_I_6 = n4_O_6; // @[Top.scala 59:10]
  assign n5_I_7 = n4_O_7; // @[Top.scala 59:10]
  assign n5_I_8 = n4_O_8; // @[Top.scala 59:10]
  assign n5_I_9 = n4_O_9; // @[Top.scala 59:10]
  assign n5_I_10 = n4_O_10; // @[Top.scala 59:10]
  assign n5_I_11 = n4_O_11; // @[Top.scala 59:10]
  assign n5_I_12 = n4_O_12; // @[Top.scala 59:10]
  assign n5_I_13 = n4_O_13; // @[Top.scala 59:10]
  assign n5_I_14 = n4_O_14; // @[Top.scala 59:10]
  assign n5_I_15 = n4_O_15; // @[Top.scala 59:10]
  assign n6_clock = clock;
  assign n6_reset = reset;
  assign n6_valid_up = n4_valid_down; // @[Top.scala 63:17]
  assign n6_I_0 = n4_O_0; // @[Top.scala 62:10]
  assign n6_I_1 = n4_O_1; // @[Top.scala 62:10]
  assign n6_I_2 = n4_O_2; // @[Top.scala 62:10]
  assign n6_I_3 = n4_O_3; // @[Top.scala 62:10]
  assign n6_I_4 = n4_O_4; // @[Top.scala 62:10]
  assign n6_I_5 = n4_O_5; // @[Top.scala 62:10]
  assign n6_I_6 = n4_O_6; // @[Top.scala 62:10]
  assign n6_I_7 = n4_O_7; // @[Top.scala 62:10]
  assign n6_I_8 = n4_O_8; // @[Top.scala 62:10]
  assign n6_I_9 = n4_O_9; // @[Top.scala 62:10]
  assign n6_I_10 = n4_O_10; // @[Top.scala 62:10]
  assign n6_I_11 = n4_O_11; // @[Top.scala 62:10]
  assign n6_I_12 = n4_O_12; // @[Top.scala 62:10]
  assign n6_I_13 = n4_O_13; // @[Top.scala 62:10]
  assign n6_I_14 = n4_O_14; // @[Top.scala 62:10]
  assign n6_I_15 = n4_O_15; // @[Top.scala 62:10]
  assign n7_valid_up = n5_valid_down & n6_valid_down; // @[Top.scala 67:17]
  assign n7_I0_0 = n5_O_0; // @[Top.scala 65:11]
  assign n7_I0_1 = n5_O_1; // @[Top.scala 65:11]
  assign n7_I0_2 = n5_O_2; // @[Top.scala 65:11]
  assign n7_I0_3 = n5_O_3; // @[Top.scala 65:11]
  assign n7_I0_4 = n5_O_4; // @[Top.scala 65:11]
  assign n7_I0_5 = n5_O_5; // @[Top.scala 65:11]
  assign n7_I0_6 = n5_O_6; // @[Top.scala 65:11]
  assign n7_I0_7 = n5_O_7; // @[Top.scala 65:11]
  assign n7_I0_8 = n5_O_8; // @[Top.scala 65:11]
  assign n7_I0_9 = n5_O_9; // @[Top.scala 65:11]
  assign n7_I0_10 = n5_O_10; // @[Top.scala 65:11]
  assign n7_I0_11 = n5_O_11; // @[Top.scala 65:11]
  assign n7_I0_12 = n5_O_12; // @[Top.scala 65:11]
  assign n7_I0_13 = n5_O_13; // @[Top.scala 65:11]
  assign n7_I0_14 = n5_O_14; // @[Top.scala 65:11]
  assign n7_I0_15 = n5_O_15; // @[Top.scala 65:11]
  assign n7_I1_0 = n6_O_0; // @[Top.scala 66:11]
  assign n7_I1_1 = n6_O_1; // @[Top.scala 66:11]
  assign n7_I1_2 = n6_O_2; // @[Top.scala 66:11]
  assign n7_I1_3 = n6_O_3; // @[Top.scala 66:11]
  assign n7_I1_4 = n6_O_4; // @[Top.scala 66:11]
  assign n7_I1_5 = n6_O_5; // @[Top.scala 66:11]
  assign n7_I1_6 = n6_O_6; // @[Top.scala 66:11]
  assign n7_I1_7 = n6_O_7; // @[Top.scala 66:11]
  assign n7_I1_8 = n6_O_8; // @[Top.scala 66:11]
  assign n7_I1_9 = n6_O_9; // @[Top.scala 66:11]
  assign n7_I1_10 = n6_O_10; // @[Top.scala 66:11]
  assign n7_I1_11 = n6_O_11; // @[Top.scala 66:11]
  assign n7_I1_12 = n6_O_12; // @[Top.scala 66:11]
  assign n7_I1_13 = n6_O_13; // @[Top.scala 66:11]
  assign n7_I1_14 = n6_O_14; // @[Top.scala 66:11]
  assign n7_I1_15 = n6_O_15; // @[Top.scala 66:11]
  assign n14_clock = clock;
  assign n14_reset = reset;
  assign n14_valid_up = n3_valid_down; // @[Top.scala 70:18]
  assign n14_I_0 = n3_O_0; // @[Top.scala 69:11]
  assign n14_I_1 = n3_O_1; // @[Top.scala 69:11]
  assign n14_I_2 = n3_O_2; // @[Top.scala 69:11]
  assign n14_I_3 = n3_O_3; // @[Top.scala 69:11]
  assign n14_I_4 = n3_O_4; // @[Top.scala 69:11]
  assign n14_I_5 = n3_O_5; // @[Top.scala 69:11]
  assign n14_I_6 = n3_O_6; // @[Top.scala 69:11]
  assign n14_I_7 = n3_O_7; // @[Top.scala 69:11]
  assign n14_I_8 = n3_O_8; // @[Top.scala 69:11]
  assign n14_I_9 = n3_O_9; // @[Top.scala 69:11]
  assign n14_I_10 = n3_O_10; // @[Top.scala 69:11]
  assign n14_I_11 = n3_O_11; // @[Top.scala 69:11]
  assign n14_I_12 = n3_O_12; // @[Top.scala 69:11]
  assign n14_I_13 = n3_O_13; // @[Top.scala 69:11]
  assign n14_I_14 = n3_O_14; // @[Top.scala 69:11]
  assign n14_I_15 = n3_O_15; // @[Top.scala 69:11]
  assign n15_valid_up = n7_valid_down & n14_valid_down; // @[Top.scala 74:18]
  assign n15_I0_0_0 = n7_O_0_0; // @[Top.scala 72:12]
  assign n15_I0_0_1 = n7_O_0_1; // @[Top.scala 72:12]
  assign n15_I0_1_0 = n7_O_1_0; // @[Top.scala 72:12]
  assign n15_I0_1_1 = n7_O_1_1; // @[Top.scala 72:12]
  assign n15_I0_2_0 = n7_O_2_0; // @[Top.scala 72:12]
  assign n15_I0_2_1 = n7_O_2_1; // @[Top.scala 72:12]
  assign n15_I0_3_0 = n7_O_3_0; // @[Top.scala 72:12]
  assign n15_I0_3_1 = n7_O_3_1; // @[Top.scala 72:12]
  assign n15_I0_4_0 = n7_O_4_0; // @[Top.scala 72:12]
  assign n15_I0_4_1 = n7_O_4_1; // @[Top.scala 72:12]
  assign n15_I0_5_0 = n7_O_5_0; // @[Top.scala 72:12]
  assign n15_I0_5_1 = n7_O_5_1; // @[Top.scala 72:12]
  assign n15_I0_6_0 = n7_O_6_0; // @[Top.scala 72:12]
  assign n15_I0_6_1 = n7_O_6_1; // @[Top.scala 72:12]
  assign n15_I0_7_0 = n7_O_7_0; // @[Top.scala 72:12]
  assign n15_I0_7_1 = n7_O_7_1; // @[Top.scala 72:12]
  assign n15_I0_8_0 = n7_O_8_0; // @[Top.scala 72:12]
  assign n15_I0_8_1 = n7_O_8_1; // @[Top.scala 72:12]
  assign n15_I0_9_0 = n7_O_9_0; // @[Top.scala 72:12]
  assign n15_I0_9_1 = n7_O_9_1; // @[Top.scala 72:12]
  assign n15_I0_10_0 = n7_O_10_0; // @[Top.scala 72:12]
  assign n15_I0_10_1 = n7_O_10_1; // @[Top.scala 72:12]
  assign n15_I0_11_0 = n7_O_11_0; // @[Top.scala 72:12]
  assign n15_I0_11_1 = n7_O_11_1; // @[Top.scala 72:12]
  assign n15_I0_12_0 = n7_O_12_0; // @[Top.scala 72:12]
  assign n15_I0_12_1 = n7_O_12_1; // @[Top.scala 72:12]
  assign n15_I0_13_0 = n7_O_13_0; // @[Top.scala 72:12]
  assign n15_I0_13_1 = n7_O_13_1; // @[Top.scala 72:12]
  assign n15_I0_14_0 = n7_O_14_0; // @[Top.scala 72:12]
  assign n15_I0_14_1 = n7_O_14_1; // @[Top.scala 72:12]
  assign n15_I0_15_0 = n7_O_15_0; // @[Top.scala 72:12]
  assign n15_I0_15_1 = n7_O_15_1; // @[Top.scala 72:12]
  assign n15_I1_0 = n14_O_0; // @[Top.scala 73:12]
  assign n15_I1_1 = n14_O_1; // @[Top.scala 73:12]
  assign n15_I1_2 = n14_O_2; // @[Top.scala 73:12]
  assign n15_I1_3 = n14_O_3; // @[Top.scala 73:12]
  assign n15_I1_4 = n14_O_4; // @[Top.scala 73:12]
  assign n15_I1_5 = n14_O_5; // @[Top.scala 73:12]
  assign n15_I1_6 = n14_O_6; // @[Top.scala 73:12]
  assign n15_I1_7 = n14_O_7; // @[Top.scala 73:12]
  assign n15_I1_8 = n14_O_8; // @[Top.scala 73:12]
  assign n15_I1_9 = n14_O_9; // @[Top.scala 73:12]
  assign n15_I1_10 = n14_O_10; // @[Top.scala 73:12]
  assign n15_I1_11 = n14_O_11; // @[Top.scala 73:12]
  assign n15_I1_12 = n14_O_12; // @[Top.scala 73:12]
  assign n15_I1_13 = n14_O_13; // @[Top.scala 73:12]
  assign n15_I1_14 = n14_O_14; // @[Top.scala 73:12]
  assign n15_I1_15 = n14_O_15; // @[Top.scala 73:12]
  assign n24_valid_up = n15_valid_down; // @[Top.scala 77:18]
  assign n24_I_0_0 = n15_O_0_0; // @[Top.scala 76:11]
  assign n24_I_0_1 = n15_O_0_1; // @[Top.scala 76:11]
  assign n24_I_0_2 = n15_O_0_2; // @[Top.scala 76:11]
  assign n24_I_1_0 = n15_O_1_0; // @[Top.scala 76:11]
  assign n24_I_1_1 = n15_O_1_1; // @[Top.scala 76:11]
  assign n24_I_1_2 = n15_O_1_2; // @[Top.scala 76:11]
  assign n24_I_2_0 = n15_O_2_0; // @[Top.scala 76:11]
  assign n24_I_2_1 = n15_O_2_1; // @[Top.scala 76:11]
  assign n24_I_2_2 = n15_O_2_2; // @[Top.scala 76:11]
  assign n24_I_3_0 = n15_O_3_0; // @[Top.scala 76:11]
  assign n24_I_3_1 = n15_O_3_1; // @[Top.scala 76:11]
  assign n24_I_3_2 = n15_O_3_2; // @[Top.scala 76:11]
  assign n24_I_4_0 = n15_O_4_0; // @[Top.scala 76:11]
  assign n24_I_4_1 = n15_O_4_1; // @[Top.scala 76:11]
  assign n24_I_4_2 = n15_O_4_2; // @[Top.scala 76:11]
  assign n24_I_5_0 = n15_O_5_0; // @[Top.scala 76:11]
  assign n24_I_5_1 = n15_O_5_1; // @[Top.scala 76:11]
  assign n24_I_5_2 = n15_O_5_2; // @[Top.scala 76:11]
  assign n24_I_6_0 = n15_O_6_0; // @[Top.scala 76:11]
  assign n24_I_6_1 = n15_O_6_1; // @[Top.scala 76:11]
  assign n24_I_6_2 = n15_O_6_2; // @[Top.scala 76:11]
  assign n24_I_7_0 = n15_O_7_0; // @[Top.scala 76:11]
  assign n24_I_7_1 = n15_O_7_1; // @[Top.scala 76:11]
  assign n24_I_7_2 = n15_O_7_2; // @[Top.scala 76:11]
  assign n24_I_8_0 = n15_O_8_0; // @[Top.scala 76:11]
  assign n24_I_8_1 = n15_O_8_1; // @[Top.scala 76:11]
  assign n24_I_8_2 = n15_O_8_2; // @[Top.scala 76:11]
  assign n24_I_9_0 = n15_O_9_0; // @[Top.scala 76:11]
  assign n24_I_9_1 = n15_O_9_1; // @[Top.scala 76:11]
  assign n24_I_9_2 = n15_O_9_2; // @[Top.scala 76:11]
  assign n24_I_10_0 = n15_O_10_0; // @[Top.scala 76:11]
  assign n24_I_10_1 = n15_O_10_1; // @[Top.scala 76:11]
  assign n24_I_10_2 = n15_O_10_2; // @[Top.scala 76:11]
  assign n24_I_11_0 = n15_O_11_0; // @[Top.scala 76:11]
  assign n24_I_11_1 = n15_O_11_1; // @[Top.scala 76:11]
  assign n24_I_11_2 = n15_O_11_2; // @[Top.scala 76:11]
  assign n24_I_12_0 = n15_O_12_0; // @[Top.scala 76:11]
  assign n24_I_12_1 = n15_O_12_1; // @[Top.scala 76:11]
  assign n24_I_12_2 = n15_O_12_2; // @[Top.scala 76:11]
  assign n24_I_13_0 = n15_O_13_0; // @[Top.scala 76:11]
  assign n24_I_13_1 = n15_O_13_1; // @[Top.scala 76:11]
  assign n24_I_13_2 = n15_O_13_2; // @[Top.scala 76:11]
  assign n24_I_14_0 = n15_O_14_0; // @[Top.scala 76:11]
  assign n24_I_14_1 = n15_O_14_1; // @[Top.scala 76:11]
  assign n24_I_14_2 = n15_O_14_2; // @[Top.scala 76:11]
  assign n24_I_15_0 = n15_O_15_0; // @[Top.scala 76:11]
  assign n24_I_15_1 = n15_O_15_1; // @[Top.scala 76:11]
  assign n24_I_15_2 = n15_O_15_2; // @[Top.scala 76:11]
  assign n31_valid_up = n24_valid_down; // @[Top.scala 80:18]
  assign n31_I_0_0_0 = n24_O_0_0_0; // @[Top.scala 79:11]
  assign n31_I_0_0_1 = n24_O_0_0_1; // @[Top.scala 79:11]
  assign n31_I_0_0_2 = n24_O_0_0_2; // @[Top.scala 79:11]
  assign n31_I_1_0_0 = n24_O_1_0_0; // @[Top.scala 79:11]
  assign n31_I_1_0_1 = n24_O_1_0_1; // @[Top.scala 79:11]
  assign n31_I_1_0_2 = n24_O_1_0_2; // @[Top.scala 79:11]
  assign n31_I_2_0_0 = n24_O_2_0_0; // @[Top.scala 79:11]
  assign n31_I_2_0_1 = n24_O_2_0_1; // @[Top.scala 79:11]
  assign n31_I_2_0_2 = n24_O_2_0_2; // @[Top.scala 79:11]
  assign n31_I_3_0_0 = n24_O_3_0_0; // @[Top.scala 79:11]
  assign n31_I_3_0_1 = n24_O_3_0_1; // @[Top.scala 79:11]
  assign n31_I_3_0_2 = n24_O_3_0_2; // @[Top.scala 79:11]
  assign n31_I_4_0_0 = n24_O_4_0_0; // @[Top.scala 79:11]
  assign n31_I_4_0_1 = n24_O_4_0_1; // @[Top.scala 79:11]
  assign n31_I_4_0_2 = n24_O_4_0_2; // @[Top.scala 79:11]
  assign n31_I_5_0_0 = n24_O_5_0_0; // @[Top.scala 79:11]
  assign n31_I_5_0_1 = n24_O_5_0_1; // @[Top.scala 79:11]
  assign n31_I_5_0_2 = n24_O_5_0_2; // @[Top.scala 79:11]
  assign n31_I_6_0_0 = n24_O_6_0_0; // @[Top.scala 79:11]
  assign n31_I_6_0_1 = n24_O_6_0_1; // @[Top.scala 79:11]
  assign n31_I_6_0_2 = n24_O_6_0_2; // @[Top.scala 79:11]
  assign n31_I_7_0_0 = n24_O_7_0_0; // @[Top.scala 79:11]
  assign n31_I_7_0_1 = n24_O_7_0_1; // @[Top.scala 79:11]
  assign n31_I_7_0_2 = n24_O_7_0_2; // @[Top.scala 79:11]
  assign n31_I_8_0_0 = n24_O_8_0_0; // @[Top.scala 79:11]
  assign n31_I_8_0_1 = n24_O_8_0_1; // @[Top.scala 79:11]
  assign n31_I_8_0_2 = n24_O_8_0_2; // @[Top.scala 79:11]
  assign n31_I_9_0_0 = n24_O_9_0_0; // @[Top.scala 79:11]
  assign n31_I_9_0_1 = n24_O_9_0_1; // @[Top.scala 79:11]
  assign n31_I_9_0_2 = n24_O_9_0_2; // @[Top.scala 79:11]
  assign n31_I_10_0_0 = n24_O_10_0_0; // @[Top.scala 79:11]
  assign n31_I_10_0_1 = n24_O_10_0_1; // @[Top.scala 79:11]
  assign n31_I_10_0_2 = n24_O_10_0_2; // @[Top.scala 79:11]
  assign n31_I_11_0_0 = n24_O_11_0_0; // @[Top.scala 79:11]
  assign n31_I_11_0_1 = n24_O_11_0_1; // @[Top.scala 79:11]
  assign n31_I_11_0_2 = n24_O_11_0_2; // @[Top.scala 79:11]
  assign n31_I_12_0_0 = n24_O_12_0_0; // @[Top.scala 79:11]
  assign n31_I_12_0_1 = n24_O_12_0_1; // @[Top.scala 79:11]
  assign n31_I_12_0_2 = n24_O_12_0_2; // @[Top.scala 79:11]
  assign n31_I_13_0_0 = n24_O_13_0_0; // @[Top.scala 79:11]
  assign n31_I_13_0_1 = n24_O_13_0_1; // @[Top.scala 79:11]
  assign n31_I_13_0_2 = n24_O_13_0_2; // @[Top.scala 79:11]
  assign n31_I_14_0_0 = n24_O_14_0_0; // @[Top.scala 79:11]
  assign n31_I_14_0_1 = n24_O_14_0_1; // @[Top.scala 79:11]
  assign n31_I_14_0_2 = n24_O_14_0_2; // @[Top.scala 79:11]
  assign n31_I_15_0_0 = n24_O_15_0_0; // @[Top.scala 79:11]
  assign n31_I_15_0_1 = n24_O_15_0_1; // @[Top.scala 79:11]
  assign n31_I_15_0_2 = n24_O_15_0_2; // @[Top.scala 79:11]
  assign n32_clock = clock;
  assign n32_reset = reset;
  assign n32_valid_up = n2_valid_down; // @[Top.scala 83:18]
  assign n32_I_0 = n2_O_0; // @[Top.scala 82:11]
  assign n32_I_1 = n2_O_1; // @[Top.scala 82:11]
  assign n32_I_2 = n2_O_2; // @[Top.scala 82:11]
  assign n32_I_3 = n2_O_3; // @[Top.scala 82:11]
  assign n32_I_4 = n2_O_4; // @[Top.scala 82:11]
  assign n32_I_5 = n2_O_5; // @[Top.scala 82:11]
  assign n32_I_6 = n2_O_6; // @[Top.scala 82:11]
  assign n32_I_7 = n2_O_7; // @[Top.scala 82:11]
  assign n32_I_8 = n2_O_8; // @[Top.scala 82:11]
  assign n32_I_9 = n2_O_9; // @[Top.scala 82:11]
  assign n32_I_10 = n2_O_10; // @[Top.scala 82:11]
  assign n32_I_11 = n2_O_11; // @[Top.scala 82:11]
  assign n32_I_12 = n2_O_12; // @[Top.scala 82:11]
  assign n32_I_13 = n2_O_13; // @[Top.scala 82:11]
  assign n32_I_14 = n2_O_14; // @[Top.scala 82:11]
  assign n32_I_15 = n2_O_15; // @[Top.scala 82:11]
  assign n33_clock = clock;
  assign n33_reset = reset;
  assign n33_valid_up = n32_valid_down; // @[Top.scala 86:18]
  assign n33_I_0 = n32_O_0; // @[Top.scala 85:11]
  assign n33_I_1 = n32_O_1; // @[Top.scala 85:11]
  assign n33_I_2 = n32_O_2; // @[Top.scala 85:11]
  assign n33_I_3 = n32_O_3; // @[Top.scala 85:11]
  assign n33_I_4 = n32_O_4; // @[Top.scala 85:11]
  assign n33_I_5 = n32_O_5; // @[Top.scala 85:11]
  assign n33_I_6 = n32_O_6; // @[Top.scala 85:11]
  assign n33_I_7 = n32_O_7; // @[Top.scala 85:11]
  assign n33_I_8 = n32_O_8; // @[Top.scala 85:11]
  assign n33_I_9 = n32_O_9; // @[Top.scala 85:11]
  assign n33_I_10 = n32_O_10; // @[Top.scala 85:11]
  assign n33_I_11 = n32_O_11; // @[Top.scala 85:11]
  assign n33_I_12 = n32_O_12; // @[Top.scala 85:11]
  assign n33_I_13 = n32_O_13; // @[Top.scala 85:11]
  assign n33_I_14 = n32_O_14; // @[Top.scala 85:11]
  assign n33_I_15 = n32_O_15; // @[Top.scala 85:11]
  assign n34_clock = clock;
  assign n34_reset = reset;
  assign n34_valid_up = n32_valid_down; // @[Top.scala 89:18]
  assign n34_I_0 = n32_O_0; // @[Top.scala 88:11]
  assign n34_I_1 = n32_O_1; // @[Top.scala 88:11]
  assign n34_I_2 = n32_O_2; // @[Top.scala 88:11]
  assign n34_I_3 = n32_O_3; // @[Top.scala 88:11]
  assign n34_I_4 = n32_O_4; // @[Top.scala 88:11]
  assign n34_I_5 = n32_O_5; // @[Top.scala 88:11]
  assign n34_I_6 = n32_O_6; // @[Top.scala 88:11]
  assign n34_I_7 = n32_O_7; // @[Top.scala 88:11]
  assign n34_I_8 = n32_O_8; // @[Top.scala 88:11]
  assign n34_I_9 = n32_O_9; // @[Top.scala 88:11]
  assign n34_I_10 = n32_O_10; // @[Top.scala 88:11]
  assign n34_I_11 = n32_O_11; // @[Top.scala 88:11]
  assign n34_I_12 = n32_O_12; // @[Top.scala 88:11]
  assign n34_I_13 = n32_O_13; // @[Top.scala 88:11]
  assign n34_I_14 = n32_O_14; // @[Top.scala 88:11]
  assign n34_I_15 = n32_O_15; // @[Top.scala 88:11]
  assign n35_valid_up = n33_valid_down & n34_valid_down; // @[Top.scala 93:18]
  assign n35_I0_0 = n33_O_0; // @[Top.scala 91:12]
  assign n35_I0_1 = n33_O_1; // @[Top.scala 91:12]
  assign n35_I0_2 = n33_O_2; // @[Top.scala 91:12]
  assign n35_I0_3 = n33_O_3; // @[Top.scala 91:12]
  assign n35_I0_4 = n33_O_4; // @[Top.scala 91:12]
  assign n35_I0_5 = n33_O_5; // @[Top.scala 91:12]
  assign n35_I0_6 = n33_O_6; // @[Top.scala 91:12]
  assign n35_I0_7 = n33_O_7; // @[Top.scala 91:12]
  assign n35_I0_8 = n33_O_8; // @[Top.scala 91:12]
  assign n35_I0_9 = n33_O_9; // @[Top.scala 91:12]
  assign n35_I0_10 = n33_O_10; // @[Top.scala 91:12]
  assign n35_I0_11 = n33_O_11; // @[Top.scala 91:12]
  assign n35_I0_12 = n33_O_12; // @[Top.scala 91:12]
  assign n35_I0_13 = n33_O_13; // @[Top.scala 91:12]
  assign n35_I0_14 = n33_O_14; // @[Top.scala 91:12]
  assign n35_I0_15 = n33_O_15; // @[Top.scala 91:12]
  assign n35_I1_0 = n34_O_0; // @[Top.scala 92:12]
  assign n35_I1_1 = n34_O_1; // @[Top.scala 92:12]
  assign n35_I1_2 = n34_O_2; // @[Top.scala 92:12]
  assign n35_I1_3 = n34_O_3; // @[Top.scala 92:12]
  assign n35_I1_4 = n34_O_4; // @[Top.scala 92:12]
  assign n35_I1_5 = n34_O_5; // @[Top.scala 92:12]
  assign n35_I1_6 = n34_O_6; // @[Top.scala 92:12]
  assign n35_I1_7 = n34_O_7; // @[Top.scala 92:12]
  assign n35_I1_8 = n34_O_8; // @[Top.scala 92:12]
  assign n35_I1_9 = n34_O_9; // @[Top.scala 92:12]
  assign n35_I1_10 = n34_O_10; // @[Top.scala 92:12]
  assign n35_I1_11 = n34_O_11; // @[Top.scala 92:12]
  assign n35_I1_12 = n34_O_12; // @[Top.scala 92:12]
  assign n35_I1_13 = n34_O_13; // @[Top.scala 92:12]
  assign n35_I1_14 = n34_O_14; // @[Top.scala 92:12]
  assign n35_I1_15 = n34_O_15; // @[Top.scala 92:12]
  assign n42_clock = clock;
  assign n42_reset = reset;
  assign n42_valid_up = n2_valid_down; // @[Top.scala 96:18]
  assign n42_I_0 = n2_O_0; // @[Top.scala 95:11]
  assign n42_I_1 = n2_O_1; // @[Top.scala 95:11]
  assign n42_I_2 = n2_O_2; // @[Top.scala 95:11]
  assign n42_I_3 = n2_O_3; // @[Top.scala 95:11]
  assign n42_I_4 = n2_O_4; // @[Top.scala 95:11]
  assign n42_I_5 = n2_O_5; // @[Top.scala 95:11]
  assign n42_I_6 = n2_O_6; // @[Top.scala 95:11]
  assign n42_I_7 = n2_O_7; // @[Top.scala 95:11]
  assign n42_I_8 = n2_O_8; // @[Top.scala 95:11]
  assign n42_I_9 = n2_O_9; // @[Top.scala 95:11]
  assign n42_I_10 = n2_O_10; // @[Top.scala 95:11]
  assign n42_I_11 = n2_O_11; // @[Top.scala 95:11]
  assign n42_I_12 = n2_O_12; // @[Top.scala 95:11]
  assign n42_I_13 = n2_O_13; // @[Top.scala 95:11]
  assign n42_I_14 = n2_O_14; // @[Top.scala 95:11]
  assign n42_I_15 = n2_O_15; // @[Top.scala 95:11]
  assign n43_valid_up = n35_valid_down & n42_valid_down; // @[Top.scala 100:18]
  assign n43_I0_0_0 = n35_O_0_0; // @[Top.scala 98:12]
  assign n43_I0_0_1 = n35_O_0_1; // @[Top.scala 98:12]
  assign n43_I0_1_0 = n35_O_1_0; // @[Top.scala 98:12]
  assign n43_I0_1_1 = n35_O_1_1; // @[Top.scala 98:12]
  assign n43_I0_2_0 = n35_O_2_0; // @[Top.scala 98:12]
  assign n43_I0_2_1 = n35_O_2_1; // @[Top.scala 98:12]
  assign n43_I0_3_0 = n35_O_3_0; // @[Top.scala 98:12]
  assign n43_I0_3_1 = n35_O_3_1; // @[Top.scala 98:12]
  assign n43_I0_4_0 = n35_O_4_0; // @[Top.scala 98:12]
  assign n43_I0_4_1 = n35_O_4_1; // @[Top.scala 98:12]
  assign n43_I0_5_0 = n35_O_5_0; // @[Top.scala 98:12]
  assign n43_I0_5_1 = n35_O_5_1; // @[Top.scala 98:12]
  assign n43_I0_6_0 = n35_O_6_0; // @[Top.scala 98:12]
  assign n43_I0_6_1 = n35_O_6_1; // @[Top.scala 98:12]
  assign n43_I0_7_0 = n35_O_7_0; // @[Top.scala 98:12]
  assign n43_I0_7_1 = n35_O_7_1; // @[Top.scala 98:12]
  assign n43_I0_8_0 = n35_O_8_0; // @[Top.scala 98:12]
  assign n43_I0_8_1 = n35_O_8_1; // @[Top.scala 98:12]
  assign n43_I0_9_0 = n35_O_9_0; // @[Top.scala 98:12]
  assign n43_I0_9_1 = n35_O_9_1; // @[Top.scala 98:12]
  assign n43_I0_10_0 = n35_O_10_0; // @[Top.scala 98:12]
  assign n43_I0_10_1 = n35_O_10_1; // @[Top.scala 98:12]
  assign n43_I0_11_0 = n35_O_11_0; // @[Top.scala 98:12]
  assign n43_I0_11_1 = n35_O_11_1; // @[Top.scala 98:12]
  assign n43_I0_12_0 = n35_O_12_0; // @[Top.scala 98:12]
  assign n43_I0_12_1 = n35_O_12_1; // @[Top.scala 98:12]
  assign n43_I0_13_0 = n35_O_13_0; // @[Top.scala 98:12]
  assign n43_I0_13_1 = n35_O_13_1; // @[Top.scala 98:12]
  assign n43_I0_14_0 = n35_O_14_0; // @[Top.scala 98:12]
  assign n43_I0_14_1 = n35_O_14_1; // @[Top.scala 98:12]
  assign n43_I0_15_0 = n35_O_15_0; // @[Top.scala 98:12]
  assign n43_I0_15_1 = n35_O_15_1; // @[Top.scala 98:12]
  assign n43_I1_0 = n42_O_0; // @[Top.scala 99:12]
  assign n43_I1_1 = n42_O_1; // @[Top.scala 99:12]
  assign n43_I1_2 = n42_O_2; // @[Top.scala 99:12]
  assign n43_I1_3 = n42_O_3; // @[Top.scala 99:12]
  assign n43_I1_4 = n42_O_4; // @[Top.scala 99:12]
  assign n43_I1_5 = n42_O_5; // @[Top.scala 99:12]
  assign n43_I1_6 = n42_O_6; // @[Top.scala 99:12]
  assign n43_I1_7 = n42_O_7; // @[Top.scala 99:12]
  assign n43_I1_8 = n42_O_8; // @[Top.scala 99:12]
  assign n43_I1_9 = n42_O_9; // @[Top.scala 99:12]
  assign n43_I1_10 = n42_O_10; // @[Top.scala 99:12]
  assign n43_I1_11 = n42_O_11; // @[Top.scala 99:12]
  assign n43_I1_12 = n42_O_12; // @[Top.scala 99:12]
  assign n43_I1_13 = n42_O_13; // @[Top.scala 99:12]
  assign n43_I1_14 = n42_O_14; // @[Top.scala 99:12]
  assign n43_I1_15 = n42_O_15; // @[Top.scala 99:12]
  assign n52_valid_up = n43_valid_down; // @[Top.scala 103:18]
  assign n52_I_0_0 = n43_O_0_0; // @[Top.scala 102:11]
  assign n52_I_0_1 = n43_O_0_1; // @[Top.scala 102:11]
  assign n52_I_0_2 = n43_O_0_2; // @[Top.scala 102:11]
  assign n52_I_1_0 = n43_O_1_0; // @[Top.scala 102:11]
  assign n52_I_1_1 = n43_O_1_1; // @[Top.scala 102:11]
  assign n52_I_1_2 = n43_O_1_2; // @[Top.scala 102:11]
  assign n52_I_2_0 = n43_O_2_0; // @[Top.scala 102:11]
  assign n52_I_2_1 = n43_O_2_1; // @[Top.scala 102:11]
  assign n52_I_2_2 = n43_O_2_2; // @[Top.scala 102:11]
  assign n52_I_3_0 = n43_O_3_0; // @[Top.scala 102:11]
  assign n52_I_3_1 = n43_O_3_1; // @[Top.scala 102:11]
  assign n52_I_3_2 = n43_O_3_2; // @[Top.scala 102:11]
  assign n52_I_4_0 = n43_O_4_0; // @[Top.scala 102:11]
  assign n52_I_4_1 = n43_O_4_1; // @[Top.scala 102:11]
  assign n52_I_4_2 = n43_O_4_2; // @[Top.scala 102:11]
  assign n52_I_5_0 = n43_O_5_0; // @[Top.scala 102:11]
  assign n52_I_5_1 = n43_O_5_1; // @[Top.scala 102:11]
  assign n52_I_5_2 = n43_O_5_2; // @[Top.scala 102:11]
  assign n52_I_6_0 = n43_O_6_0; // @[Top.scala 102:11]
  assign n52_I_6_1 = n43_O_6_1; // @[Top.scala 102:11]
  assign n52_I_6_2 = n43_O_6_2; // @[Top.scala 102:11]
  assign n52_I_7_0 = n43_O_7_0; // @[Top.scala 102:11]
  assign n52_I_7_1 = n43_O_7_1; // @[Top.scala 102:11]
  assign n52_I_7_2 = n43_O_7_2; // @[Top.scala 102:11]
  assign n52_I_8_0 = n43_O_8_0; // @[Top.scala 102:11]
  assign n52_I_8_1 = n43_O_8_1; // @[Top.scala 102:11]
  assign n52_I_8_2 = n43_O_8_2; // @[Top.scala 102:11]
  assign n52_I_9_0 = n43_O_9_0; // @[Top.scala 102:11]
  assign n52_I_9_1 = n43_O_9_1; // @[Top.scala 102:11]
  assign n52_I_9_2 = n43_O_9_2; // @[Top.scala 102:11]
  assign n52_I_10_0 = n43_O_10_0; // @[Top.scala 102:11]
  assign n52_I_10_1 = n43_O_10_1; // @[Top.scala 102:11]
  assign n52_I_10_2 = n43_O_10_2; // @[Top.scala 102:11]
  assign n52_I_11_0 = n43_O_11_0; // @[Top.scala 102:11]
  assign n52_I_11_1 = n43_O_11_1; // @[Top.scala 102:11]
  assign n52_I_11_2 = n43_O_11_2; // @[Top.scala 102:11]
  assign n52_I_12_0 = n43_O_12_0; // @[Top.scala 102:11]
  assign n52_I_12_1 = n43_O_12_1; // @[Top.scala 102:11]
  assign n52_I_12_2 = n43_O_12_2; // @[Top.scala 102:11]
  assign n52_I_13_0 = n43_O_13_0; // @[Top.scala 102:11]
  assign n52_I_13_1 = n43_O_13_1; // @[Top.scala 102:11]
  assign n52_I_13_2 = n43_O_13_2; // @[Top.scala 102:11]
  assign n52_I_14_0 = n43_O_14_0; // @[Top.scala 102:11]
  assign n52_I_14_1 = n43_O_14_1; // @[Top.scala 102:11]
  assign n52_I_14_2 = n43_O_14_2; // @[Top.scala 102:11]
  assign n52_I_15_0 = n43_O_15_0; // @[Top.scala 102:11]
  assign n52_I_15_1 = n43_O_15_1; // @[Top.scala 102:11]
  assign n52_I_15_2 = n43_O_15_2; // @[Top.scala 102:11]
  assign n59_valid_up = n52_valid_down; // @[Top.scala 106:18]
  assign n59_I_0_0_0 = n52_O_0_0_0; // @[Top.scala 105:11]
  assign n59_I_0_0_1 = n52_O_0_0_1; // @[Top.scala 105:11]
  assign n59_I_0_0_2 = n52_O_0_0_2; // @[Top.scala 105:11]
  assign n59_I_1_0_0 = n52_O_1_0_0; // @[Top.scala 105:11]
  assign n59_I_1_0_1 = n52_O_1_0_1; // @[Top.scala 105:11]
  assign n59_I_1_0_2 = n52_O_1_0_2; // @[Top.scala 105:11]
  assign n59_I_2_0_0 = n52_O_2_0_0; // @[Top.scala 105:11]
  assign n59_I_2_0_1 = n52_O_2_0_1; // @[Top.scala 105:11]
  assign n59_I_2_0_2 = n52_O_2_0_2; // @[Top.scala 105:11]
  assign n59_I_3_0_0 = n52_O_3_0_0; // @[Top.scala 105:11]
  assign n59_I_3_0_1 = n52_O_3_0_1; // @[Top.scala 105:11]
  assign n59_I_3_0_2 = n52_O_3_0_2; // @[Top.scala 105:11]
  assign n59_I_4_0_0 = n52_O_4_0_0; // @[Top.scala 105:11]
  assign n59_I_4_0_1 = n52_O_4_0_1; // @[Top.scala 105:11]
  assign n59_I_4_0_2 = n52_O_4_0_2; // @[Top.scala 105:11]
  assign n59_I_5_0_0 = n52_O_5_0_0; // @[Top.scala 105:11]
  assign n59_I_5_0_1 = n52_O_5_0_1; // @[Top.scala 105:11]
  assign n59_I_5_0_2 = n52_O_5_0_2; // @[Top.scala 105:11]
  assign n59_I_6_0_0 = n52_O_6_0_0; // @[Top.scala 105:11]
  assign n59_I_6_0_1 = n52_O_6_0_1; // @[Top.scala 105:11]
  assign n59_I_6_0_2 = n52_O_6_0_2; // @[Top.scala 105:11]
  assign n59_I_7_0_0 = n52_O_7_0_0; // @[Top.scala 105:11]
  assign n59_I_7_0_1 = n52_O_7_0_1; // @[Top.scala 105:11]
  assign n59_I_7_0_2 = n52_O_7_0_2; // @[Top.scala 105:11]
  assign n59_I_8_0_0 = n52_O_8_0_0; // @[Top.scala 105:11]
  assign n59_I_8_0_1 = n52_O_8_0_1; // @[Top.scala 105:11]
  assign n59_I_8_0_2 = n52_O_8_0_2; // @[Top.scala 105:11]
  assign n59_I_9_0_0 = n52_O_9_0_0; // @[Top.scala 105:11]
  assign n59_I_9_0_1 = n52_O_9_0_1; // @[Top.scala 105:11]
  assign n59_I_9_0_2 = n52_O_9_0_2; // @[Top.scala 105:11]
  assign n59_I_10_0_0 = n52_O_10_0_0; // @[Top.scala 105:11]
  assign n59_I_10_0_1 = n52_O_10_0_1; // @[Top.scala 105:11]
  assign n59_I_10_0_2 = n52_O_10_0_2; // @[Top.scala 105:11]
  assign n59_I_11_0_0 = n52_O_11_0_0; // @[Top.scala 105:11]
  assign n59_I_11_0_1 = n52_O_11_0_1; // @[Top.scala 105:11]
  assign n59_I_11_0_2 = n52_O_11_0_2; // @[Top.scala 105:11]
  assign n59_I_12_0_0 = n52_O_12_0_0; // @[Top.scala 105:11]
  assign n59_I_12_0_1 = n52_O_12_0_1; // @[Top.scala 105:11]
  assign n59_I_12_0_2 = n52_O_12_0_2; // @[Top.scala 105:11]
  assign n59_I_13_0_0 = n52_O_13_0_0; // @[Top.scala 105:11]
  assign n59_I_13_0_1 = n52_O_13_0_1; // @[Top.scala 105:11]
  assign n59_I_13_0_2 = n52_O_13_0_2; // @[Top.scala 105:11]
  assign n59_I_14_0_0 = n52_O_14_0_0; // @[Top.scala 105:11]
  assign n59_I_14_0_1 = n52_O_14_0_1; // @[Top.scala 105:11]
  assign n59_I_14_0_2 = n52_O_14_0_2; // @[Top.scala 105:11]
  assign n59_I_15_0_0 = n52_O_15_0_0; // @[Top.scala 105:11]
  assign n59_I_15_0_1 = n52_O_15_0_1; // @[Top.scala 105:11]
  assign n59_I_15_0_2 = n52_O_15_0_2; // @[Top.scala 105:11]
  assign n60_clock = clock;
  assign n60_reset = reset;
  assign n60_valid_up = n59_valid_down; // @[Top.scala 109:18]
  assign n60_I_0_0 = n59_O_0_0; // @[Top.scala 108:11]
  assign n60_I_0_1 = n59_O_0_1; // @[Top.scala 108:11]
  assign n60_I_0_2 = n59_O_0_2; // @[Top.scala 108:11]
  assign n60_I_1_0 = n59_O_1_0; // @[Top.scala 108:11]
  assign n60_I_1_1 = n59_O_1_1; // @[Top.scala 108:11]
  assign n60_I_1_2 = n59_O_1_2; // @[Top.scala 108:11]
  assign n60_I_2_0 = n59_O_2_0; // @[Top.scala 108:11]
  assign n60_I_2_1 = n59_O_2_1; // @[Top.scala 108:11]
  assign n60_I_2_2 = n59_O_2_2; // @[Top.scala 108:11]
  assign n60_I_3_0 = n59_O_3_0; // @[Top.scala 108:11]
  assign n60_I_3_1 = n59_O_3_1; // @[Top.scala 108:11]
  assign n60_I_3_2 = n59_O_3_2; // @[Top.scala 108:11]
  assign n60_I_4_0 = n59_O_4_0; // @[Top.scala 108:11]
  assign n60_I_4_1 = n59_O_4_1; // @[Top.scala 108:11]
  assign n60_I_4_2 = n59_O_4_2; // @[Top.scala 108:11]
  assign n60_I_5_0 = n59_O_5_0; // @[Top.scala 108:11]
  assign n60_I_5_1 = n59_O_5_1; // @[Top.scala 108:11]
  assign n60_I_5_2 = n59_O_5_2; // @[Top.scala 108:11]
  assign n60_I_6_0 = n59_O_6_0; // @[Top.scala 108:11]
  assign n60_I_6_1 = n59_O_6_1; // @[Top.scala 108:11]
  assign n60_I_6_2 = n59_O_6_2; // @[Top.scala 108:11]
  assign n60_I_7_0 = n59_O_7_0; // @[Top.scala 108:11]
  assign n60_I_7_1 = n59_O_7_1; // @[Top.scala 108:11]
  assign n60_I_7_2 = n59_O_7_2; // @[Top.scala 108:11]
  assign n60_I_8_0 = n59_O_8_0; // @[Top.scala 108:11]
  assign n60_I_8_1 = n59_O_8_1; // @[Top.scala 108:11]
  assign n60_I_8_2 = n59_O_8_2; // @[Top.scala 108:11]
  assign n60_I_9_0 = n59_O_9_0; // @[Top.scala 108:11]
  assign n60_I_9_1 = n59_O_9_1; // @[Top.scala 108:11]
  assign n60_I_9_2 = n59_O_9_2; // @[Top.scala 108:11]
  assign n60_I_10_0 = n59_O_10_0; // @[Top.scala 108:11]
  assign n60_I_10_1 = n59_O_10_1; // @[Top.scala 108:11]
  assign n60_I_10_2 = n59_O_10_2; // @[Top.scala 108:11]
  assign n60_I_11_0 = n59_O_11_0; // @[Top.scala 108:11]
  assign n60_I_11_1 = n59_O_11_1; // @[Top.scala 108:11]
  assign n60_I_11_2 = n59_O_11_2; // @[Top.scala 108:11]
  assign n60_I_12_0 = n59_O_12_0; // @[Top.scala 108:11]
  assign n60_I_12_1 = n59_O_12_1; // @[Top.scala 108:11]
  assign n60_I_12_2 = n59_O_12_2; // @[Top.scala 108:11]
  assign n60_I_13_0 = n59_O_13_0; // @[Top.scala 108:11]
  assign n60_I_13_1 = n59_O_13_1; // @[Top.scala 108:11]
  assign n60_I_13_2 = n59_O_13_2; // @[Top.scala 108:11]
  assign n60_I_14_0 = n59_O_14_0; // @[Top.scala 108:11]
  assign n60_I_14_1 = n59_O_14_1; // @[Top.scala 108:11]
  assign n60_I_14_2 = n59_O_14_2; // @[Top.scala 108:11]
  assign n60_I_15_0 = n59_O_15_0; // @[Top.scala 108:11]
  assign n60_I_15_1 = n59_O_15_1; // @[Top.scala 108:11]
  assign n60_I_15_2 = n59_O_15_2; // @[Top.scala 108:11]
  assign n61_valid_up = n31_valid_down & n60_valid_down; // @[Top.scala 113:18]
  assign n61_I0_0_0 = n31_O_0_0; // @[Top.scala 111:12]
  assign n61_I0_0_1 = n31_O_0_1; // @[Top.scala 111:12]
  assign n61_I0_0_2 = n31_O_0_2; // @[Top.scala 111:12]
  assign n61_I0_1_0 = n31_O_1_0; // @[Top.scala 111:12]
  assign n61_I0_1_1 = n31_O_1_1; // @[Top.scala 111:12]
  assign n61_I0_1_2 = n31_O_1_2; // @[Top.scala 111:12]
  assign n61_I0_2_0 = n31_O_2_0; // @[Top.scala 111:12]
  assign n61_I0_2_1 = n31_O_2_1; // @[Top.scala 111:12]
  assign n61_I0_2_2 = n31_O_2_2; // @[Top.scala 111:12]
  assign n61_I0_3_0 = n31_O_3_0; // @[Top.scala 111:12]
  assign n61_I0_3_1 = n31_O_3_1; // @[Top.scala 111:12]
  assign n61_I0_3_2 = n31_O_3_2; // @[Top.scala 111:12]
  assign n61_I0_4_0 = n31_O_4_0; // @[Top.scala 111:12]
  assign n61_I0_4_1 = n31_O_4_1; // @[Top.scala 111:12]
  assign n61_I0_4_2 = n31_O_4_2; // @[Top.scala 111:12]
  assign n61_I0_5_0 = n31_O_5_0; // @[Top.scala 111:12]
  assign n61_I0_5_1 = n31_O_5_1; // @[Top.scala 111:12]
  assign n61_I0_5_2 = n31_O_5_2; // @[Top.scala 111:12]
  assign n61_I0_6_0 = n31_O_6_0; // @[Top.scala 111:12]
  assign n61_I0_6_1 = n31_O_6_1; // @[Top.scala 111:12]
  assign n61_I0_6_2 = n31_O_6_2; // @[Top.scala 111:12]
  assign n61_I0_7_0 = n31_O_7_0; // @[Top.scala 111:12]
  assign n61_I0_7_1 = n31_O_7_1; // @[Top.scala 111:12]
  assign n61_I0_7_2 = n31_O_7_2; // @[Top.scala 111:12]
  assign n61_I0_8_0 = n31_O_8_0; // @[Top.scala 111:12]
  assign n61_I0_8_1 = n31_O_8_1; // @[Top.scala 111:12]
  assign n61_I0_8_2 = n31_O_8_2; // @[Top.scala 111:12]
  assign n61_I0_9_0 = n31_O_9_0; // @[Top.scala 111:12]
  assign n61_I0_9_1 = n31_O_9_1; // @[Top.scala 111:12]
  assign n61_I0_9_2 = n31_O_9_2; // @[Top.scala 111:12]
  assign n61_I0_10_0 = n31_O_10_0; // @[Top.scala 111:12]
  assign n61_I0_10_1 = n31_O_10_1; // @[Top.scala 111:12]
  assign n61_I0_10_2 = n31_O_10_2; // @[Top.scala 111:12]
  assign n61_I0_11_0 = n31_O_11_0; // @[Top.scala 111:12]
  assign n61_I0_11_1 = n31_O_11_1; // @[Top.scala 111:12]
  assign n61_I0_11_2 = n31_O_11_2; // @[Top.scala 111:12]
  assign n61_I0_12_0 = n31_O_12_0; // @[Top.scala 111:12]
  assign n61_I0_12_1 = n31_O_12_1; // @[Top.scala 111:12]
  assign n61_I0_12_2 = n31_O_12_2; // @[Top.scala 111:12]
  assign n61_I0_13_0 = n31_O_13_0; // @[Top.scala 111:12]
  assign n61_I0_13_1 = n31_O_13_1; // @[Top.scala 111:12]
  assign n61_I0_13_2 = n31_O_13_2; // @[Top.scala 111:12]
  assign n61_I0_14_0 = n31_O_14_0; // @[Top.scala 111:12]
  assign n61_I0_14_1 = n31_O_14_1; // @[Top.scala 111:12]
  assign n61_I0_14_2 = n31_O_14_2; // @[Top.scala 111:12]
  assign n61_I0_15_0 = n31_O_15_0; // @[Top.scala 111:12]
  assign n61_I0_15_1 = n31_O_15_1; // @[Top.scala 111:12]
  assign n61_I0_15_2 = n31_O_15_2; // @[Top.scala 111:12]
  assign n61_I1_0_0 = n60_O_0_0; // @[Top.scala 112:12]
  assign n61_I1_0_1 = n60_O_0_1; // @[Top.scala 112:12]
  assign n61_I1_0_2 = n60_O_0_2; // @[Top.scala 112:12]
  assign n61_I1_1_0 = n60_O_1_0; // @[Top.scala 112:12]
  assign n61_I1_1_1 = n60_O_1_1; // @[Top.scala 112:12]
  assign n61_I1_1_2 = n60_O_1_2; // @[Top.scala 112:12]
  assign n61_I1_2_0 = n60_O_2_0; // @[Top.scala 112:12]
  assign n61_I1_2_1 = n60_O_2_1; // @[Top.scala 112:12]
  assign n61_I1_2_2 = n60_O_2_2; // @[Top.scala 112:12]
  assign n61_I1_3_0 = n60_O_3_0; // @[Top.scala 112:12]
  assign n61_I1_3_1 = n60_O_3_1; // @[Top.scala 112:12]
  assign n61_I1_3_2 = n60_O_3_2; // @[Top.scala 112:12]
  assign n61_I1_4_0 = n60_O_4_0; // @[Top.scala 112:12]
  assign n61_I1_4_1 = n60_O_4_1; // @[Top.scala 112:12]
  assign n61_I1_4_2 = n60_O_4_2; // @[Top.scala 112:12]
  assign n61_I1_5_0 = n60_O_5_0; // @[Top.scala 112:12]
  assign n61_I1_5_1 = n60_O_5_1; // @[Top.scala 112:12]
  assign n61_I1_5_2 = n60_O_5_2; // @[Top.scala 112:12]
  assign n61_I1_6_0 = n60_O_6_0; // @[Top.scala 112:12]
  assign n61_I1_6_1 = n60_O_6_1; // @[Top.scala 112:12]
  assign n61_I1_6_2 = n60_O_6_2; // @[Top.scala 112:12]
  assign n61_I1_7_0 = n60_O_7_0; // @[Top.scala 112:12]
  assign n61_I1_7_1 = n60_O_7_1; // @[Top.scala 112:12]
  assign n61_I1_7_2 = n60_O_7_2; // @[Top.scala 112:12]
  assign n61_I1_8_0 = n60_O_8_0; // @[Top.scala 112:12]
  assign n61_I1_8_1 = n60_O_8_1; // @[Top.scala 112:12]
  assign n61_I1_8_2 = n60_O_8_2; // @[Top.scala 112:12]
  assign n61_I1_9_0 = n60_O_9_0; // @[Top.scala 112:12]
  assign n61_I1_9_1 = n60_O_9_1; // @[Top.scala 112:12]
  assign n61_I1_9_2 = n60_O_9_2; // @[Top.scala 112:12]
  assign n61_I1_10_0 = n60_O_10_0; // @[Top.scala 112:12]
  assign n61_I1_10_1 = n60_O_10_1; // @[Top.scala 112:12]
  assign n61_I1_10_2 = n60_O_10_2; // @[Top.scala 112:12]
  assign n61_I1_11_0 = n60_O_11_0; // @[Top.scala 112:12]
  assign n61_I1_11_1 = n60_O_11_1; // @[Top.scala 112:12]
  assign n61_I1_11_2 = n60_O_11_2; // @[Top.scala 112:12]
  assign n61_I1_12_0 = n60_O_12_0; // @[Top.scala 112:12]
  assign n61_I1_12_1 = n60_O_12_1; // @[Top.scala 112:12]
  assign n61_I1_12_2 = n60_O_12_2; // @[Top.scala 112:12]
  assign n61_I1_13_0 = n60_O_13_0; // @[Top.scala 112:12]
  assign n61_I1_13_1 = n60_O_13_1; // @[Top.scala 112:12]
  assign n61_I1_13_2 = n60_O_13_2; // @[Top.scala 112:12]
  assign n61_I1_14_0 = n60_O_14_0; // @[Top.scala 112:12]
  assign n61_I1_14_1 = n60_O_14_1; // @[Top.scala 112:12]
  assign n61_I1_14_2 = n60_O_14_2; // @[Top.scala 112:12]
  assign n61_I1_15_0 = n60_O_15_0; // @[Top.scala 112:12]
  assign n61_I1_15_1 = n60_O_15_1; // @[Top.scala 112:12]
  assign n61_I1_15_2 = n60_O_15_2; // @[Top.scala 112:12]
  assign n68_clock = clock;
  assign n68_reset = reset;
  assign n68_valid_up = n1_valid_down; // @[Top.scala 116:18]
  assign n68_I_0 = n1_O_0; // @[Top.scala 115:11]
  assign n68_I_1 = n1_O_1; // @[Top.scala 115:11]
  assign n68_I_2 = n1_O_2; // @[Top.scala 115:11]
  assign n68_I_3 = n1_O_3; // @[Top.scala 115:11]
  assign n68_I_4 = n1_O_4; // @[Top.scala 115:11]
  assign n68_I_5 = n1_O_5; // @[Top.scala 115:11]
  assign n68_I_6 = n1_O_6; // @[Top.scala 115:11]
  assign n68_I_7 = n1_O_7; // @[Top.scala 115:11]
  assign n68_I_8 = n1_O_8; // @[Top.scala 115:11]
  assign n68_I_9 = n1_O_9; // @[Top.scala 115:11]
  assign n68_I_10 = n1_O_10; // @[Top.scala 115:11]
  assign n68_I_11 = n1_O_11; // @[Top.scala 115:11]
  assign n68_I_12 = n1_O_12; // @[Top.scala 115:11]
  assign n68_I_13 = n1_O_13; // @[Top.scala 115:11]
  assign n68_I_14 = n1_O_14; // @[Top.scala 115:11]
  assign n68_I_15 = n1_O_15; // @[Top.scala 115:11]
  assign n69_clock = clock;
  assign n69_reset = reset;
  assign n69_valid_up = n68_valid_down; // @[Top.scala 119:18]
  assign n69_I_0 = n68_O_0; // @[Top.scala 118:11]
  assign n69_I_1 = n68_O_1; // @[Top.scala 118:11]
  assign n69_I_2 = n68_O_2; // @[Top.scala 118:11]
  assign n69_I_3 = n68_O_3; // @[Top.scala 118:11]
  assign n69_I_4 = n68_O_4; // @[Top.scala 118:11]
  assign n69_I_5 = n68_O_5; // @[Top.scala 118:11]
  assign n69_I_6 = n68_O_6; // @[Top.scala 118:11]
  assign n69_I_7 = n68_O_7; // @[Top.scala 118:11]
  assign n69_I_8 = n68_O_8; // @[Top.scala 118:11]
  assign n69_I_9 = n68_O_9; // @[Top.scala 118:11]
  assign n69_I_10 = n68_O_10; // @[Top.scala 118:11]
  assign n69_I_11 = n68_O_11; // @[Top.scala 118:11]
  assign n69_I_12 = n68_O_12; // @[Top.scala 118:11]
  assign n69_I_13 = n68_O_13; // @[Top.scala 118:11]
  assign n69_I_14 = n68_O_14; // @[Top.scala 118:11]
  assign n69_I_15 = n68_O_15; // @[Top.scala 118:11]
  assign n70_clock = clock;
  assign n70_reset = reset;
  assign n70_valid_up = n68_valid_down; // @[Top.scala 122:18]
  assign n70_I_0 = n68_O_0; // @[Top.scala 121:11]
  assign n70_I_1 = n68_O_1; // @[Top.scala 121:11]
  assign n70_I_2 = n68_O_2; // @[Top.scala 121:11]
  assign n70_I_3 = n68_O_3; // @[Top.scala 121:11]
  assign n70_I_4 = n68_O_4; // @[Top.scala 121:11]
  assign n70_I_5 = n68_O_5; // @[Top.scala 121:11]
  assign n70_I_6 = n68_O_6; // @[Top.scala 121:11]
  assign n70_I_7 = n68_O_7; // @[Top.scala 121:11]
  assign n70_I_8 = n68_O_8; // @[Top.scala 121:11]
  assign n70_I_9 = n68_O_9; // @[Top.scala 121:11]
  assign n70_I_10 = n68_O_10; // @[Top.scala 121:11]
  assign n70_I_11 = n68_O_11; // @[Top.scala 121:11]
  assign n70_I_12 = n68_O_12; // @[Top.scala 121:11]
  assign n70_I_13 = n68_O_13; // @[Top.scala 121:11]
  assign n70_I_14 = n68_O_14; // @[Top.scala 121:11]
  assign n70_I_15 = n68_O_15; // @[Top.scala 121:11]
  assign n71_valid_up = n69_valid_down & n70_valid_down; // @[Top.scala 126:18]
  assign n71_I0_0 = n69_O_0; // @[Top.scala 124:12]
  assign n71_I0_1 = n69_O_1; // @[Top.scala 124:12]
  assign n71_I0_2 = n69_O_2; // @[Top.scala 124:12]
  assign n71_I0_3 = n69_O_3; // @[Top.scala 124:12]
  assign n71_I0_4 = n69_O_4; // @[Top.scala 124:12]
  assign n71_I0_5 = n69_O_5; // @[Top.scala 124:12]
  assign n71_I0_6 = n69_O_6; // @[Top.scala 124:12]
  assign n71_I0_7 = n69_O_7; // @[Top.scala 124:12]
  assign n71_I0_8 = n69_O_8; // @[Top.scala 124:12]
  assign n71_I0_9 = n69_O_9; // @[Top.scala 124:12]
  assign n71_I0_10 = n69_O_10; // @[Top.scala 124:12]
  assign n71_I0_11 = n69_O_11; // @[Top.scala 124:12]
  assign n71_I0_12 = n69_O_12; // @[Top.scala 124:12]
  assign n71_I0_13 = n69_O_13; // @[Top.scala 124:12]
  assign n71_I0_14 = n69_O_14; // @[Top.scala 124:12]
  assign n71_I0_15 = n69_O_15; // @[Top.scala 124:12]
  assign n71_I1_0 = n70_O_0; // @[Top.scala 125:12]
  assign n71_I1_1 = n70_O_1; // @[Top.scala 125:12]
  assign n71_I1_2 = n70_O_2; // @[Top.scala 125:12]
  assign n71_I1_3 = n70_O_3; // @[Top.scala 125:12]
  assign n71_I1_4 = n70_O_4; // @[Top.scala 125:12]
  assign n71_I1_5 = n70_O_5; // @[Top.scala 125:12]
  assign n71_I1_6 = n70_O_6; // @[Top.scala 125:12]
  assign n71_I1_7 = n70_O_7; // @[Top.scala 125:12]
  assign n71_I1_8 = n70_O_8; // @[Top.scala 125:12]
  assign n71_I1_9 = n70_O_9; // @[Top.scala 125:12]
  assign n71_I1_10 = n70_O_10; // @[Top.scala 125:12]
  assign n71_I1_11 = n70_O_11; // @[Top.scala 125:12]
  assign n71_I1_12 = n70_O_12; // @[Top.scala 125:12]
  assign n71_I1_13 = n70_O_13; // @[Top.scala 125:12]
  assign n71_I1_14 = n70_O_14; // @[Top.scala 125:12]
  assign n71_I1_15 = n70_O_15; // @[Top.scala 125:12]
  assign n78_clock = clock;
  assign n78_reset = reset;
  assign n78_valid_up = n1_valid_down; // @[Top.scala 129:18]
  assign n78_I_0 = n1_O_0; // @[Top.scala 128:11]
  assign n78_I_1 = n1_O_1; // @[Top.scala 128:11]
  assign n78_I_2 = n1_O_2; // @[Top.scala 128:11]
  assign n78_I_3 = n1_O_3; // @[Top.scala 128:11]
  assign n78_I_4 = n1_O_4; // @[Top.scala 128:11]
  assign n78_I_5 = n1_O_5; // @[Top.scala 128:11]
  assign n78_I_6 = n1_O_6; // @[Top.scala 128:11]
  assign n78_I_7 = n1_O_7; // @[Top.scala 128:11]
  assign n78_I_8 = n1_O_8; // @[Top.scala 128:11]
  assign n78_I_9 = n1_O_9; // @[Top.scala 128:11]
  assign n78_I_10 = n1_O_10; // @[Top.scala 128:11]
  assign n78_I_11 = n1_O_11; // @[Top.scala 128:11]
  assign n78_I_12 = n1_O_12; // @[Top.scala 128:11]
  assign n78_I_13 = n1_O_13; // @[Top.scala 128:11]
  assign n78_I_14 = n1_O_14; // @[Top.scala 128:11]
  assign n78_I_15 = n1_O_15; // @[Top.scala 128:11]
  assign n79_valid_up = n71_valid_down & n78_valid_down; // @[Top.scala 133:18]
  assign n79_I0_0_0 = n71_O_0_0; // @[Top.scala 131:12]
  assign n79_I0_0_1 = n71_O_0_1; // @[Top.scala 131:12]
  assign n79_I0_1_0 = n71_O_1_0; // @[Top.scala 131:12]
  assign n79_I0_1_1 = n71_O_1_1; // @[Top.scala 131:12]
  assign n79_I0_2_0 = n71_O_2_0; // @[Top.scala 131:12]
  assign n79_I0_2_1 = n71_O_2_1; // @[Top.scala 131:12]
  assign n79_I0_3_0 = n71_O_3_0; // @[Top.scala 131:12]
  assign n79_I0_3_1 = n71_O_3_1; // @[Top.scala 131:12]
  assign n79_I0_4_0 = n71_O_4_0; // @[Top.scala 131:12]
  assign n79_I0_4_1 = n71_O_4_1; // @[Top.scala 131:12]
  assign n79_I0_5_0 = n71_O_5_0; // @[Top.scala 131:12]
  assign n79_I0_5_1 = n71_O_5_1; // @[Top.scala 131:12]
  assign n79_I0_6_0 = n71_O_6_0; // @[Top.scala 131:12]
  assign n79_I0_6_1 = n71_O_6_1; // @[Top.scala 131:12]
  assign n79_I0_7_0 = n71_O_7_0; // @[Top.scala 131:12]
  assign n79_I0_7_1 = n71_O_7_1; // @[Top.scala 131:12]
  assign n79_I0_8_0 = n71_O_8_0; // @[Top.scala 131:12]
  assign n79_I0_8_1 = n71_O_8_1; // @[Top.scala 131:12]
  assign n79_I0_9_0 = n71_O_9_0; // @[Top.scala 131:12]
  assign n79_I0_9_1 = n71_O_9_1; // @[Top.scala 131:12]
  assign n79_I0_10_0 = n71_O_10_0; // @[Top.scala 131:12]
  assign n79_I0_10_1 = n71_O_10_1; // @[Top.scala 131:12]
  assign n79_I0_11_0 = n71_O_11_0; // @[Top.scala 131:12]
  assign n79_I0_11_1 = n71_O_11_1; // @[Top.scala 131:12]
  assign n79_I0_12_0 = n71_O_12_0; // @[Top.scala 131:12]
  assign n79_I0_12_1 = n71_O_12_1; // @[Top.scala 131:12]
  assign n79_I0_13_0 = n71_O_13_0; // @[Top.scala 131:12]
  assign n79_I0_13_1 = n71_O_13_1; // @[Top.scala 131:12]
  assign n79_I0_14_0 = n71_O_14_0; // @[Top.scala 131:12]
  assign n79_I0_14_1 = n71_O_14_1; // @[Top.scala 131:12]
  assign n79_I0_15_0 = n71_O_15_0; // @[Top.scala 131:12]
  assign n79_I0_15_1 = n71_O_15_1; // @[Top.scala 131:12]
  assign n79_I1_0 = n78_O_0; // @[Top.scala 132:12]
  assign n79_I1_1 = n78_O_1; // @[Top.scala 132:12]
  assign n79_I1_2 = n78_O_2; // @[Top.scala 132:12]
  assign n79_I1_3 = n78_O_3; // @[Top.scala 132:12]
  assign n79_I1_4 = n78_O_4; // @[Top.scala 132:12]
  assign n79_I1_5 = n78_O_5; // @[Top.scala 132:12]
  assign n79_I1_6 = n78_O_6; // @[Top.scala 132:12]
  assign n79_I1_7 = n78_O_7; // @[Top.scala 132:12]
  assign n79_I1_8 = n78_O_8; // @[Top.scala 132:12]
  assign n79_I1_9 = n78_O_9; // @[Top.scala 132:12]
  assign n79_I1_10 = n78_O_10; // @[Top.scala 132:12]
  assign n79_I1_11 = n78_O_11; // @[Top.scala 132:12]
  assign n79_I1_12 = n78_O_12; // @[Top.scala 132:12]
  assign n79_I1_13 = n78_O_13; // @[Top.scala 132:12]
  assign n79_I1_14 = n78_O_14; // @[Top.scala 132:12]
  assign n79_I1_15 = n78_O_15; // @[Top.scala 132:12]
  assign n88_valid_up = n79_valid_down; // @[Top.scala 136:18]
  assign n88_I_0_0 = n79_O_0_0; // @[Top.scala 135:11]
  assign n88_I_0_1 = n79_O_0_1; // @[Top.scala 135:11]
  assign n88_I_0_2 = n79_O_0_2; // @[Top.scala 135:11]
  assign n88_I_1_0 = n79_O_1_0; // @[Top.scala 135:11]
  assign n88_I_1_1 = n79_O_1_1; // @[Top.scala 135:11]
  assign n88_I_1_2 = n79_O_1_2; // @[Top.scala 135:11]
  assign n88_I_2_0 = n79_O_2_0; // @[Top.scala 135:11]
  assign n88_I_2_1 = n79_O_2_1; // @[Top.scala 135:11]
  assign n88_I_2_2 = n79_O_2_2; // @[Top.scala 135:11]
  assign n88_I_3_0 = n79_O_3_0; // @[Top.scala 135:11]
  assign n88_I_3_1 = n79_O_3_1; // @[Top.scala 135:11]
  assign n88_I_3_2 = n79_O_3_2; // @[Top.scala 135:11]
  assign n88_I_4_0 = n79_O_4_0; // @[Top.scala 135:11]
  assign n88_I_4_1 = n79_O_4_1; // @[Top.scala 135:11]
  assign n88_I_4_2 = n79_O_4_2; // @[Top.scala 135:11]
  assign n88_I_5_0 = n79_O_5_0; // @[Top.scala 135:11]
  assign n88_I_5_1 = n79_O_5_1; // @[Top.scala 135:11]
  assign n88_I_5_2 = n79_O_5_2; // @[Top.scala 135:11]
  assign n88_I_6_0 = n79_O_6_0; // @[Top.scala 135:11]
  assign n88_I_6_1 = n79_O_6_1; // @[Top.scala 135:11]
  assign n88_I_6_2 = n79_O_6_2; // @[Top.scala 135:11]
  assign n88_I_7_0 = n79_O_7_0; // @[Top.scala 135:11]
  assign n88_I_7_1 = n79_O_7_1; // @[Top.scala 135:11]
  assign n88_I_7_2 = n79_O_7_2; // @[Top.scala 135:11]
  assign n88_I_8_0 = n79_O_8_0; // @[Top.scala 135:11]
  assign n88_I_8_1 = n79_O_8_1; // @[Top.scala 135:11]
  assign n88_I_8_2 = n79_O_8_2; // @[Top.scala 135:11]
  assign n88_I_9_0 = n79_O_9_0; // @[Top.scala 135:11]
  assign n88_I_9_1 = n79_O_9_1; // @[Top.scala 135:11]
  assign n88_I_9_2 = n79_O_9_2; // @[Top.scala 135:11]
  assign n88_I_10_0 = n79_O_10_0; // @[Top.scala 135:11]
  assign n88_I_10_1 = n79_O_10_1; // @[Top.scala 135:11]
  assign n88_I_10_2 = n79_O_10_2; // @[Top.scala 135:11]
  assign n88_I_11_0 = n79_O_11_0; // @[Top.scala 135:11]
  assign n88_I_11_1 = n79_O_11_1; // @[Top.scala 135:11]
  assign n88_I_11_2 = n79_O_11_2; // @[Top.scala 135:11]
  assign n88_I_12_0 = n79_O_12_0; // @[Top.scala 135:11]
  assign n88_I_12_1 = n79_O_12_1; // @[Top.scala 135:11]
  assign n88_I_12_2 = n79_O_12_2; // @[Top.scala 135:11]
  assign n88_I_13_0 = n79_O_13_0; // @[Top.scala 135:11]
  assign n88_I_13_1 = n79_O_13_1; // @[Top.scala 135:11]
  assign n88_I_13_2 = n79_O_13_2; // @[Top.scala 135:11]
  assign n88_I_14_0 = n79_O_14_0; // @[Top.scala 135:11]
  assign n88_I_14_1 = n79_O_14_1; // @[Top.scala 135:11]
  assign n88_I_14_2 = n79_O_14_2; // @[Top.scala 135:11]
  assign n88_I_15_0 = n79_O_15_0; // @[Top.scala 135:11]
  assign n88_I_15_1 = n79_O_15_1; // @[Top.scala 135:11]
  assign n88_I_15_2 = n79_O_15_2; // @[Top.scala 135:11]
  assign n95_valid_up = n88_valid_down; // @[Top.scala 139:18]
  assign n95_I_0_0_0 = n88_O_0_0_0; // @[Top.scala 138:11]
  assign n95_I_0_0_1 = n88_O_0_0_1; // @[Top.scala 138:11]
  assign n95_I_0_0_2 = n88_O_0_0_2; // @[Top.scala 138:11]
  assign n95_I_1_0_0 = n88_O_1_0_0; // @[Top.scala 138:11]
  assign n95_I_1_0_1 = n88_O_1_0_1; // @[Top.scala 138:11]
  assign n95_I_1_0_2 = n88_O_1_0_2; // @[Top.scala 138:11]
  assign n95_I_2_0_0 = n88_O_2_0_0; // @[Top.scala 138:11]
  assign n95_I_2_0_1 = n88_O_2_0_1; // @[Top.scala 138:11]
  assign n95_I_2_0_2 = n88_O_2_0_2; // @[Top.scala 138:11]
  assign n95_I_3_0_0 = n88_O_3_0_0; // @[Top.scala 138:11]
  assign n95_I_3_0_1 = n88_O_3_0_1; // @[Top.scala 138:11]
  assign n95_I_3_0_2 = n88_O_3_0_2; // @[Top.scala 138:11]
  assign n95_I_4_0_0 = n88_O_4_0_0; // @[Top.scala 138:11]
  assign n95_I_4_0_1 = n88_O_4_0_1; // @[Top.scala 138:11]
  assign n95_I_4_0_2 = n88_O_4_0_2; // @[Top.scala 138:11]
  assign n95_I_5_0_0 = n88_O_5_0_0; // @[Top.scala 138:11]
  assign n95_I_5_0_1 = n88_O_5_0_1; // @[Top.scala 138:11]
  assign n95_I_5_0_2 = n88_O_5_0_2; // @[Top.scala 138:11]
  assign n95_I_6_0_0 = n88_O_6_0_0; // @[Top.scala 138:11]
  assign n95_I_6_0_1 = n88_O_6_0_1; // @[Top.scala 138:11]
  assign n95_I_6_0_2 = n88_O_6_0_2; // @[Top.scala 138:11]
  assign n95_I_7_0_0 = n88_O_7_0_0; // @[Top.scala 138:11]
  assign n95_I_7_0_1 = n88_O_7_0_1; // @[Top.scala 138:11]
  assign n95_I_7_0_2 = n88_O_7_0_2; // @[Top.scala 138:11]
  assign n95_I_8_0_0 = n88_O_8_0_0; // @[Top.scala 138:11]
  assign n95_I_8_0_1 = n88_O_8_0_1; // @[Top.scala 138:11]
  assign n95_I_8_0_2 = n88_O_8_0_2; // @[Top.scala 138:11]
  assign n95_I_9_0_0 = n88_O_9_0_0; // @[Top.scala 138:11]
  assign n95_I_9_0_1 = n88_O_9_0_1; // @[Top.scala 138:11]
  assign n95_I_9_0_2 = n88_O_9_0_2; // @[Top.scala 138:11]
  assign n95_I_10_0_0 = n88_O_10_0_0; // @[Top.scala 138:11]
  assign n95_I_10_0_1 = n88_O_10_0_1; // @[Top.scala 138:11]
  assign n95_I_10_0_2 = n88_O_10_0_2; // @[Top.scala 138:11]
  assign n95_I_11_0_0 = n88_O_11_0_0; // @[Top.scala 138:11]
  assign n95_I_11_0_1 = n88_O_11_0_1; // @[Top.scala 138:11]
  assign n95_I_11_0_2 = n88_O_11_0_2; // @[Top.scala 138:11]
  assign n95_I_12_0_0 = n88_O_12_0_0; // @[Top.scala 138:11]
  assign n95_I_12_0_1 = n88_O_12_0_1; // @[Top.scala 138:11]
  assign n95_I_12_0_2 = n88_O_12_0_2; // @[Top.scala 138:11]
  assign n95_I_13_0_0 = n88_O_13_0_0; // @[Top.scala 138:11]
  assign n95_I_13_0_1 = n88_O_13_0_1; // @[Top.scala 138:11]
  assign n95_I_13_0_2 = n88_O_13_0_2; // @[Top.scala 138:11]
  assign n95_I_14_0_0 = n88_O_14_0_0; // @[Top.scala 138:11]
  assign n95_I_14_0_1 = n88_O_14_0_1; // @[Top.scala 138:11]
  assign n95_I_14_0_2 = n88_O_14_0_2; // @[Top.scala 138:11]
  assign n95_I_15_0_0 = n88_O_15_0_0; // @[Top.scala 138:11]
  assign n95_I_15_0_1 = n88_O_15_0_1; // @[Top.scala 138:11]
  assign n95_I_15_0_2 = n88_O_15_0_2; // @[Top.scala 138:11]
  assign n96_clock = clock;
  assign n96_reset = reset;
  assign n96_valid_up = n95_valid_down; // @[Top.scala 142:18]
  assign n96_I_0_0 = n95_O_0_0; // @[Top.scala 141:11]
  assign n96_I_0_1 = n95_O_0_1; // @[Top.scala 141:11]
  assign n96_I_0_2 = n95_O_0_2; // @[Top.scala 141:11]
  assign n96_I_1_0 = n95_O_1_0; // @[Top.scala 141:11]
  assign n96_I_1_1 = n95_O_1_1; // @[Top.scala 141:11]
  assign n96_I_1_2 = n95_O_1_2; // @[Top.scala 141:11]
  assign n96_I_2_0 = n95_O_2_0; // @[Top.scala 141:11]
  assign n96_I_2_1 = n95_O_2_1; // @[Top.scala 141:11]
  assign n96_I_2_2 = n95_O_2_2; // @[Top.scala 141:11]
  assign n96_I_3_0 = n95_O_3_0; // @[Top.scala 141:11]
  assign n96_I_3_1 = n95_O_3_1; // @[Top.scala 141:11]
  assign n96_I_3_2 = n95_O_3_2; // @[Top.scala 141:11]
  assign n96_I_4_0 = n95_O_4_0; // @[Top.scala 141:11]
  assign n96_I_4_1 = n95_O_4_1; // @[Top.scala 141:11]
  assign n96_I_4_2 = n95_O_4_2; // @[Top.scala 141:11]
  assign n96_I_5_0 = n95_O_5_0; // @[Top.scala 141:11]
  assign n96_I_5_1 = n95_O_5_1; // @[Top.scala 141:11]
  assign n96_I_5_2 = n95_O_5_2; // @[Top.scala 141:11]
  assign n96_I_6_0 = n95_O_6_0; // @[Top.scala 141:11]
  assign n96_I_6_1 = n95_O_6_1; // @[Top.scala 141:11]
  assign n96_I_6_2 = n95_O_6_2; // @[Top.scala 141:11]
  assign n96_I_7_0 = n95_O_7_0; // @[Top.scala 141:11]
  assign n96_I_7_1 = n95_O_7_1; // @[Top.scala 141:11]
  assign n96_I_7_2 = n95_O_7_2; // @[Top.scala 141:11]
  assign n96_I_8_0 = n95_O_8_0; // @[Top.scala 141:11]
  assign n96_I_8_1 = n95_O_8_1; // @[Top.scala 141:11]
  assign n96_I_8_2 = n95_O_8_2; // @[Top.scala 141:11]
  assign n96_I_9_0 = n95_O_9_0; // @[Top.scala 141:11]
  assign n96_I_9_1 = n95_O_9_1; // @[Top.scala 141:11]
  assign n96_I_9_2 = n95_O_9_2; // @[Top.scala 141:11]
  assign n96_I_10_0 = n95_O_10_0; // @[Top.scala 141:11]
  assign n96_I_10_1 = n95_O_10_1; // @[Top.scala 141:11]
  assign n96_I_10_2 = n95_O_10_2; // @[Top.scala 141:11]
  assign n96_I_11_0 = n95_O_11_0; // @[Top.scala 141:11]
  assign n96_I_11_1 = n95_O_11_1; // @[Top.scala 141:11]
  assign n96_I_11_2 = n95_O_11_2; // @[Top.scala 141:11]
  assign n96_I_12_0 = n95_O_12_0; // @[Top.scala 141:11]
  assign n96_I_12_1 = n95_O_12_1; // @[Top.scala 141:11]
  assign n96_I_12_2 = n95_O_12_2; // @[Top.scala 141:11]
  assign n96_I_13_0 = n95_O_13_0; // @[Top.scala 141:11]
  assign n96_I_13_1 = n95_O_13_1; // @[Top.scala 141:11]
  assign n96_I_13_2 = n95_O_13_2; // @[Top.scala 141:11]
  assign n96_I_14_0 = n95_O_14_0; // @[Top.scala 141:11]
  assign n96_I_14_1 = n95_O_14_1; // @[Top.scala 141:11]
  assign n96_I_14_2 = n95_O_14_2; // @[Top.scala 141:11]
  assign n96_I_15_0 = n95_O_15_0; // @[Top.scala 141:11]
  assign n96_I_15_1 = n95_O_15_1; // @[Top.scala 141:11]
  assign n96_I_15_2 = n95_O_15_2; // @[Top.scala 141:11]
  assign n97_valid_up = n61_valid_down & n96_valid_down; // @[Top.scala 146:18]
  assign n97_I0_0_0_0 = n61_O_0_0_0; // @[Top.scala 144:12]
  assign n97_I0_0_0_1 = n61_O_0_0_1; // @[Top.scala 144:12]
  assign n97_I0_0_0_2 = n61_O_0_0_2; // @[Top.scala 144:12]
  assign n97_I0_0_1_0 = n61_O_0_1_0; // @[Top.scala 144:12]
  assign n97_I0_0_1_1 = n61_O_0_1_1; // @[Top.scala 144:12]
  assign n97_I0_0_1_2 = n61_O_0_1_2; // @[Top.scala 144:12]
  assign n97_I0_1_0_0 = n61_O_1_0_0; // @[Top.scala 144:12]
  assign n97_I0_1_0_1 = n61_O_1_0_1; // @[Top.scala 144:12]
  assign n97_I0_1_0_2 = n61_O_1_0_2; // @[Top.scala 144:12]
  assign n97_I0_1_1_0 = n61_O_1_1_0; // @[Top.scala 144:12]
  assign n97_I0_1_1_1 = n61_O_1_1_1; // @[Top.scala 144:12]
  assign n97_I0_1_1_2 = n61_O_1_1_2; // @[Top.scala 144:12]
  assign n97_I0_2_0_0 = n61_O_2_0_0; // @[Top.scala 144:12]
  assign n97_I0_2_0_1 = n61_O_2_0_1; // @[Top.scala 144:12]
  assign n97_I0_2_0_2 = n61_O_2_0_2; // @[Top.scala 144:12]
  assign n97_I0_2_1_0 = n61_O_2_1_0; // @[Top.scala 144:12]
  assign n97_I0_2_1_1 = n61_O_2_1_1; // @[Top.scala 144:12]
  assign n97_I0_2_1_2 = n61_O_2_1_2; // @[Top.scala 144:12]
  assign n97_I0_3_0_0 = n61_O_3_0_0; // @[Top.scala 144:12]
  assign n97_I0_3_0_1 = n61_O_3_0_1; // @[Top.scala 144:12]
  assign n97_I0_3_0_2 = n61_O_3_0_2; // @[Top.scala 144:12]
  assign n97_I0_3_1_0 = n61_O_3_1_0; // @[Top.scala 144:12]
  assign n97_I0_3_1_1 = n61_O_3_1_1; // @[Top.scala 144:12]
  assign n97_I0_3_1_2 = n61_O_3_1_2; // @[Top.scala 144:12]
  assign n97_I0_4_0_0 = n61_O_4_0_0; // @[Top.scala 144:12]
  assign n97_I0_4_0_1 = n61_O_4_0_1; // @[Top.scala 144:12]
  assign n97_I0_4_0_2 = n61_O_4_0_2; // @[Top.scala 144:12]
  assign n97_I0_4_1_0 = n61_O_4_1_0; // @[Top.scala 144:12]
  assign n97_I0_4_1_1 = n61_O_4_1_1; // @[Top.scala 144:12]
  assign n97_I0_4_1_2 = n61_O_4_1_2; // @[Top.scala 144:12]
  assign n97_I0_5_0_0 = n61_O_5_0_0; // @[Top.scala 144:12]
  assign n97_I0_5_0_1 = n61_O_5_0_1; // @[Top.scala 144:12]
  assign n97_I0_5_0_2 = n61_O_5_0_2; // @[Top.scala 144:12]
  assign n97_I0_5_1_0 = n61_O_5_1_0; // @[Top.scala 144:12]
  assign n97_I0_5_1_1 = n61_O_5_1_1; // @[Top.scala 144:12]
  assign n97_I0_5_1_2 = n61_O_5_1_2; // @[Top.scala 144:12]
  assign n97_I0_6_0_0 = n61_O_6_0_0; // @[Top.scala 144:12]
  assign n97_I0_6_0_1 = n61_O_6_0_1; // @[Top.scala 144:12]
  assign n97_I0_6_0_2 = n61_O_6_0_2; // @[Top.scala 144:12]
  assign n97_I0_6_1_0 = n61_O_6_1_0; // @[Top.scala 144:12]
  assign n97_I0_6_1_1 = n61_O_6_1_1; // @[Top.scala 144:12]
  assign n97_I0_6_1_2 = n61_O_6_1_2; // @[Top.scala 144:12]
  assign n97_I0_7_0_0 = n61_O_7_0_0; // @[Top.scala 144:12]
  assign n97_I0_7_0_1 = n61_O_7_0_1; // @[Top.scala 144:12]
  assign n97_I0_7_0_2 = n61_O_7_0_2; // @[Top.scala 144:12]
  assign n97_I0_7_1_0 = n61_O_7_1_0; // @[Top.scala 144:12]
  assign n97_I0_7_1_1 = n61_O_7_1_1; // @[Top.scala 144:12]
  assign n97_I0_7_1_2 = n61_O_7_1_2; // @[Top.scala 144:12]
  assign n97_I0_8_0_0 = n61_O_8_0_0; // @[Top.scala 144:12]
  assign n97_I0_8_0_1 = n61_O_8_0_1; // @[Top.scala 144:12]
  assign n97_I0_8_0_2 = n61_O_8_0_2; // @[Top.scala 144:12]
  assign n97_I0_8_1_0 = n61_O_8_1_0; // @[Top.scala 144:12]
  assign n97_I0_8_1_1 = n61_O_8_1_1; // @[Top.scala 144:12]
  assign n97_I0_8_1_2 = n61_O_8_1_2; // @[Top.scala 144:12]
  assign n97_I0_9_0_0 = n61_O_9_0_0; // @[Top.scala 144:12]
  assign n97_I0_9_0_1 = n61_O_9_0_1; // @[Top.scala 144:12]
  assign n97_I0_9_0_2 = n61_O_9_0_2; // @[Top.scala 144:12]
  assign n97_I0_9_1_0 = n61_O_9_1_0; // @[Top.scala 144:12]
  assign n97_I0_9_1_1 = n61_O_9_1_1; // @[Top.scala 144:12]
  assign n97_I0_9_1_2 = n61_O_9_1_2; // @[Top.scala 144:12]
  assign n97_I0_10_0_0 = n61_O_10_0_0; // @[Top.scala 144:12]
  assign n97_I0_10_0_1 = n61_O_10_0_1; // @[Top.scala 144:12]
  assign n97_I0_10_0_2 = n61_O_10_0_2; // @[Top.scala 144:12]
  assign n97_I0_10_1_0 = n61_O_10_1_0; // @[Top.scala 144:12]
  assign n97_I0_10_1_1 = n61_O_10_1_1; // @[Top.scala 144:12]
  assign n97_I0_10_1_2 = n61_O_10_1_2; // @[Top.scala 144:12]
  assign n97_I0_11_0_0 = n61_O_11_0_0; // @[Top.scala 144:12]
  assign n97_I0_11_0_1 = n61_O_11_0_1; // @[Top.scala 144:12]
  assign n97_I0_11_0_2 = n61_O_11_0_2; // @[Top.scala 144:12]
  assign n97_I0_11_1_0 = n61_O_11_1_0; // @[Top.scala 144:12]
  assign n97_I0_11_1_1 = n61_O_11_1_1; // @[Top.scala 144:12]
  assign n97_I0_11_1_2 = n61_O_11_1_2; // @[Top.scala 144:12]
  assign n97_I0_12_0_0 = n61_O_12_0_0; // @[Top.scala 144:12]
  assign n97_I0_12_0_1 = n61_O_12_0_1; // @[Top.scala 144:12]
  assign n97_I0_12_0_2 = n61_O_12_0_2; // @[Top.scala 144:12]
  assign n97_I0_12_1_0 = n61_O_12_1_0; // @[Top.scala 144:12]
  assign n97_I0_12_1_1 = n61_O_12_1_1; // @[Top.scala 144:12]
  assign n97_I0_12_1_2 = n61_O_12_1_2; // @[Top.scala 144:12]
  assign n97_I0_13_0_0 = n61_O_13_0_0; // @[Top.scala 144:12]
  assign n97_I0_13_0_1 = n61_O_13_0_1; // @[Top.scala 144:12]
  assign n97_I0_13_0_2 = n61_O_13_0_2; // @[Top.scala 144:12]
  assign n97_I0_13_1_0 = n61_O_13_1_0; // @[Top.scala 144:12]
  assign n97_I0_13_1_1 = n61_O_13_1_1; // @[Top.scala 144:12]
  assign n97_I0_13_1_2 = n61_O_13_1_2; // @[Top.scala 144:12]
  assign n97_I0_14_0_0 = n61_O_14_0_0; // @[Top.scala 144:12]
  assign n97_I0_14_0_1 = n61_O_14_0_1; // @[Top.scala 144:12]
  assign n97_I0_14_0_2 = n61_O_14_0_2; // @[Top.scala 144:12]
  assign n97_I0_14_1_0 = n61_O_14_1_0; // @[Top.scala 144:12]
  assign n97_I0_14_1_1 = n61_O_14_1_1; // @[Top.scala 144:12]
  assign n97_I0_14_1_2 = n61_O_14_1_2; // @[Top.scala 144:12]
  assign n97_I0_15_0_0 = n61_O_15_0_0; // @[Top.scala 144:12]
  assign n97_I0_15_0_1 = n61_O_15_0_1; // @[Top.scala 144:12]
  assign n97_I0_15_0_2 = n61_O_15_0_2; // @[Top.scala 144:12]
  assign n97_I0_15_1_0 = n61_O_15_1_0; // @[Top.scala 144:12]
  assign n97_I0_15_1_1 = n61_O_15_1_1; // @[Top.scala 144:12]
  assign n97_I0_15_1_2 = n61_O_15_1_2; // @[Top.scala 144:12]
  assign n97_I1_0_0 = n96_O_0_0; // @[Top.scala 145:12]
  assign n97_I1_0_1 = n96_O_0_1; // @[Top.scala 145:12]
  assign n97_I1_0_2 = n96_O_0_2; // @[Top.scala 145:12]
  assign n97_I1_1_0 = n96_O_1_0; // @[Top.scala 145:12]
  assign n97_I1_1_1 = n96_O_1_1; // @[Top.scala 145:12]
  assign n97_I1_1_2 = n96_O_1_2; // @[Top.scala 145:12]
  assign n97_I1_2_0 = n96_O_2_0; // @[Top.scala 145:12]
  assign n97_I1_2_1 = n96_O_2_1; // @[Top.scala 145:12]
  assign n97_I1_2_2 = n96_O_2_2; // @[Top.scala 145:12]
  assign n97_I1_3_0 = n96_O_3_0; // @[Top.scala 145:12]
  assign n97_I1_3_1 = n96_O_3_1; // @[Top.scala 145:12]
  assign n97_I1_3_2 = n96_O_3_2; // @[Top.scala 145:12]
  assign n97_I1_4_0 = n96_O_4_0; // @[Top.scala 145:12]
  assign n97_I1_4_1 = n96_O_4_1; // @[Top.scala 145:12]
  assign n97_I1_4_2 = n96_O_4_2; // @[Top.scala 145:12]
  assign n97_I1_5_0 = n96_O_5_0; // @[Top.scala 145:12]
  assign n97_I1_5_1 = n96_O_5_1; // @[Top.scala 145:12]
  assign n97_I1_5_2 = n96_O_5_2; // @[Top.scala 145:12]
  assign n97_I1_6_0 = n96_O_6_0; // @[Top.scala 145:12]
  assign n97_I1_6_1 = n96_O_6_1; // @[Top.scala 145:12]
  assign n97_I1_6_2 = n96_O_6_2; // @[Top.scala 145:12]
  assign n97_I1_7_0 = n96_O_7_0; // @[Top.scala 145:12]
  assign n97_I1_7_1 = n96_O_7_1; // @[Top.scala 145:12]
  assign n97_I1_7_2 = n96_O_7_2; // @[Top.scala 145:12]
  assign n97_I1_8_0 = n96_O_8_0; // @[Top.scala 145:12]
  assign n97_I1_8_1 = n96_O_8_1; // @[Top.scala 145:12]
  assign n97_I1_8_2 = n96_O_8_2; // @[Top.scala 145:12]
  assign n97_I1_9_0 = n96_O_9_0; // @[Top.scala 145:12]
  assign n97_I1_9_1 = n96_O_9_1; // @[Top.scala 145:12]
  assign n97_I1_9_2 = n96_O_9_2; // @[Top.scala 145:12]
  assign n97_I1_10_0 = n96_O_10_0; // @[Top.scala 145:12]
  assign n97_I1_10_1 = n96_O_10_1; // @[Top.scala 145:12]
  assign n97_I1_10_2 = n96_O_10_2; // @[Top.scala 145:12]
  assign n97_I1_11_0 = n96_O_11_0; // @[Top.scala 145:12]
  assign n97_I1_11_1 = n96_O_11_1; // @[Top.scala 145:12]
  assign n97_I1_11_2 = n96_O_11_2; // @[Top.scala 145:12]
  assign n97_I1_12_0 = n96_O_12_0; // @[Top.scala 145:12]
  assign n97_I1_12_1 = n96_O_12_1; // @[Top.scala 145:12]
  assign n97_I1_12_2 = n96_O_12_2; // @[Top.scala 145:12]
  assign n97_I1_13_0 = n96_O_13_0; // @[Top.scala 145:12]
  assign n97_I1_13_1 = n96_O_13_1; // @[Top.scala 145:12]
  assign n97_I1_13_2 = n96_O_13_2; // @[Top.scala 145:12]
  assign n97_I1_14_0 = n96_O_14_0; // @[Top.scala 145:12]
  assign n97_I1_14_1 = n96_O_14_1; // @[Top.scala 145:12]
  assign n97_I1_14_2 = n96_O_14_2; // @[Top.scala 145:12]
  assign n97_I1_15_0 = n96_O_15_0; // @[Top.scala 145:12]
  assign n97_I1_15_1 = n96_O_15_1; // @[Top.scala 145:12]
  assign n97_I1_15_2 = n96_O_15_2; // @[Top.scala 145:12]
  assign n106_valid_up = n97_valid_down; // @[Top.scala 149:19]
  assign n106_I_0_0_0 = n97_O_0_0_0; // @[Top.scala 148:12]
  assign n106_I_0_0_1 = n97_O_0_0_1; // @[Top.scala 148:12]
  assign n106_I_0_0_2 = n97_O_0_0_2; // @[Top.scala 148:12]
  assign n106_I_0_1_0 = n97_O_0_1_0; // @[Top.scala 148:12]
  assign n106_I_0_1_1 = n97_O_0_1_1; // @[Top.scala 148:12]
  assign n106_I_0_1_2 = n97_O_0_1_2; // @[Top.scala 148:12]
  assign n106_I_0_2_0 = n97_O_0_2_0; // @[Top.scala 148:12]
  assign n106_I_0_2_1 = n97_O_0_2_1; // @[Top.scala 148:12]
  assign n106_I_0_2_2 = n97_O_0_2_2; // @[Top.scala 148:12]
  assign n106_I_1_0_0 = n97_O_1_0_0; // @[Top.scala 148:12]
  assign n106_I_1_0_1 = n97_O_1_0_1; // @[Top.scala 148:12]
  assign n106_I_1_0_2 = n97_O_1_0_2; // @[Top.scala 148:12]
  assign n106_I_1_1_0 = n97_O_1_1_0; // @[Top.scala 148:12]
  assign n106_I_1_1_1 = n97_O_1_1_1; // @[Top.scala 148:12]
  assign n106_I_1_1_2 = n97_O_1_1_2; // @[Top.scala 148:12]
  assign n106_I_1_2_0 = n97_O_1_2_0; // @[Top.scala 148:12]
  assign n106_I_1_2_1 = n97_O_1_2_1; // @[Top.scala 148:12]
  assign n106_I_1_2_2 = n97_O_1_2_2; // @[Top.scala 148:12]
  assign n106_I_2_0_0 = n97_O_2_0_0; // @[Top.scala 148:12]
  assign n106_I_2_0_1 = n97_O_2_0_1; // @[Top.scala 148:12]
  assign n106_I_2_0_2 = n97_O_2_0_2; // @[Top.scala 148:12]
  assign n106_I_2_1_0 = n97_O_2_1_0; // @[Top.scala 148:12]
  assign n106_I_2_1_1 = n97_O_2_1_1; // @[Top.scala 148:12]
  assign n106_I_2_1_2 = n97_O_2_1_2; // @[Top.scala 148:12]
  assign n106_I_2_2_0 = n97_O_2_2_0; // @[Top.scala 148:12]
  assign n106_I_2_2_1 = n97_O_2_2_1; // @[Top.scala 148:12]
  assign n106_I_2_2_2 = n97_O_2_2_2; // @[Top.scala 148:12]
  assign n106_I_3_0_0 = n97_O_3_0_0; // @[Top.scala 148:12]
  assign n106_I_3_0_1 = n97_O_3_0_1; // @[Top.scala 148:12]
  assign n106_I_3_0_2 = n97_O_3_0_2; // @[Top.scala 148:12]
  assign n106_I_3_1_0 = n97_O_3_1_0; // @[Top.scala 148:12]
  assign n106_I_3_1_1 = n97_O_3_1_1; // @[Top.scala 148:12]
  assign n106_I_3_1_2 = n97_O_3_1_2; // @[Top.scala 148:12]
  assign n106_I_3_2_0 = n97_O_3_2_0; // @[Top.scala 148:12]
  assign n106_I_3_2_1 = n97_O_3_2_1; // @[Top.scala 148:12]
  assign n106_I_3_2_2 = n97_O_3_2_2; // @[Top.scala 148:12]
  assign n106_I_4_0_0 = n97_O_4_0_0; // @[Top.scala 148:12]
  assign n106_I_4_0_1 = n97_O_4_0_1; // @[Top.scala 148:12]
  assign n106_I_4_0_2 = n97_O_4_0_2; // @[Top.scala 148:12]
  assign n106_I_4_1_0 = n97_O_4_1_0; // @[Top.scala 148:12]
  assign n106_I_4_1_1 = n97_O_4_1_1; // @[Top.scala 148:12]
  assign n106_I_4_1_2 = n97_O_4_1_2; // @[Top.scala 148:12]
  assign n106_I_4_2_0 = n97_O_4_2_0; // @[Top.scala 148:12]
  assign n106_I_4_2_1 = n97_O_4_2_1; // @[Top.scala 148:12]
  assign n106_I_4_2_2 = n97_O_4_2_2; // @[Top.scala 148:12]
  assign n106_I_5_0_0 = n97_O_5_0_0; // @[Top.scala 148:12]
  assign n106_I_5_0_1 = n97_O_5_0_1; // @[Top.scala 148:12]
  assign n106_I_5_0_2 = n97_O_5_0_2; // @[Top.scala 148:12]
  assign n106_I_5_1_0 = n97_O_5_1_0; // @[Top.scala 148:12]
  assign n106_I_5_1_1 = n97_O_5_1_1; // @[Top.scala 148:12]
  assign n106_I_5_1_2 = n97_O_5_1_2; // @[Top.scala 148:12]
  assign n106_I_5_2_0 = n97_O_5_2_0; // @[Top.scala 148:12]
  assign n106_I_5_2_1 = n97_O_5_2_1; // @[Top.scala 148:12]
  assign n106_I_5_2_2 = n97_O_5_2_2; // @[Top.scala 148:12]
  assign n106_I_6_0_0 = n97_O_6_0_0; // @[Top.scala 148:12]
  assign n106_I_6_0_1 = n97_O_6_0_1; // @[Top.scala 148:12]
  assign n106_I_6_0_2 = n97_O_6_0_2; // @[Top.scala 148:12]
  assign n106_I_6_1_0 = n97_O_6_1_0; // @[Top.scala 148:12]
  assign n106_I_6_1_1 = n97_O_6_1_1; // @[Top.scala 148:12]
  assign n106_I_6_1_2 = n97_O_6_1_2; // @[Top.scala 148:12]
  assign n106_I_6_2_0 = n97_O_6_2_0; // @[Top.scala 148:12]
  assign n106_I_6_2_1 = n97_O_6_2_1; // @[Top.scala 148:12]
  assign n106_I_6_2_2 = n97_O_6_2_2; // @[Top.scala 148:12]
  assign n106_I_7_0_0 = n97_O_7_0_0; // @[Top.scala 148:12]
  assign n106_I_7_0_1 = n97_O_7_0_1; // @[Top.scala 148:12]
  assign n106_I_7_0_2 = n97_O_7_0_2; // @[Top.scala 148:12]
  assign n106_I_7_1_0 = n97_O_7_1_0; // @[Top.scala 148:12]
  assign n106_I_7_1_1 = n97_O_7_1_1; // @[Top.scala 148:12]
  assign n106_I_7_1_2 = n97_O_7_1_2; // @[Top.scala 148:12]
  assign n106_I_7_2_0 = n97_O_7_2_0; // @[Top.scala 148:12]
  assign n106_I_7_2_1 = n97_O_7_2_1; // @[Top.scala 148:12]
  assign n106_I_7_2_2 = n97_O_7_2_2; // @[Top.scala 148:12]
  assign n106_I_8_0_0 = n97_O_8_0_0; // @[Top.scala 148:12]
  assign n106_I_8_0_1 = n97_O_8_0_1; // @[Top.scala 148:12]
  assign n106_I_8_0_2 = n97_O_8_0_2; // @[Top.scala 148:12]
  assign n106_I_8_1_0 = n97_O_8_1_0; // @[Top.scala 148:12]
  assign n106_I_8_1_1 = n97_O_8_1_1; // @[Top.scala 148:12]
  assign n106_I_8_1_2 = n97_O_8_1_2; // @[Top.scala 148:12]
  assign n106_I_8_2_0 = n97_O_8_2_0; // @[Top.scala 148:12]
  assign n106_I_8_2_1 = n97_O_8_2_1; // @[Top.scala 148:12]
  assign n106_I_8_2_2 = n97_O_8_2_2; // @[Top.scala 148:12]
  assign n106_I_9_0_0 = n97_O_9_0_0; // @[Top.scala 148:12]
  assign n106_I_9_0_1 = n97_O_9_0_1; // @[Top.scala 148:12]
  assign n106_I_9_0_2 = n97_O_9_0_2; // @[Top.scala 148:12]
  assign n106_I_9_1_0 = n97_O_9_1_0; // @[Top.scala 148:12]
  assign n106_I_9_1_1 = n97_O_9_1_1; // @[Top.scala 148:12]
  assign n106_I_9_1_2 = n97_O_9_1_2; // @[Top.scala 148:12]
  assign n106_I_9_2_0 = n97_O_9_2_0; // @[Top.scala 148:12]
  assign n106_I_9_2_1 = n97_O_9_2_1; // @[Top.scala 148:12]
  assign n106_I_9_2_2 = n97_O_9_2_2; // @[Top.scala 148:12]
  assign n106_I_10_0_0 = n97_O_10_0_0; // @[Top.scala 148:12]
  assign n106_I_10_0_1 = n97_O_10_0_1; // @[Top.scala 148:12]
  assign n106_I_10_0_2 = n97_O_10_0_2; // @[Top.scala 148:12]
  assign n106_I_10_1_0 = n97_O_10_1_0; // @[Top.scala 148:12]
  assign n106_I_10_1_1 = n97_O_10_1_1; // @[Top.scala 148:12]
  assign n106_I_10_1_2 = n97_O_10_1_2; // @[Top.scala 148:12]
  assign n106_I_10_2_0 = n97_O_10_2_0; // @[Top.scala 148:12]
  assign n106_I_10_2_1 = n97_O_10_2_1; // @[Top.scala 148:12]
  assign n106_I_10_2_2 = n97_O_10_2_2; // @[Top.scala 148:12]
  assign n106_I_11_0_0 = n97_O_11_0_0; // @[Top.scala 148:12]
  assign n106_I_11_0_1 = n97_O_11_0_1; // @[Top.scala 148:12]
  assign n106_I_11_0_2 = n97_O_11_0_2; // @[Top.scala 148:12]
  assign n106_I_11_1_0 = n97_O_11_1_0; // @[Top.scala 148:12]
  assign n106_I_11_1_1 = n97_O_11_1_1; // @[Top.scala 148:12]
  assign n106_I_11_1_2 = n97_O_11_1_2; // @[Top.scala 148:12]
  assign n106_I_11_2_0 = n97_O_11_2_0; // @[Top.scala 148:12]
  assign n106_I_11_2_1 = n97_O_11_2_1; // @[Top.scala 148:12]
  assign n106_I_11_2_2 = n97_O_11_2_2; // @[Top.scala 148:12]
  assign n106_I_12_0_0 = n97_O_12_0_0; // @[Top.scala 148:12]
  assign n106_I_12_0_1 = n97_O_12_0_1; // @[Top.scala 148:12]
  assign n106_I_12_0_2 = n97_O_12_0_2; // @[Top.scala 148:12]
  assign n106_I_12_1_0 = n97_O_12_1_0; // @[Top.scala 148:12]
  assign n106_I_12_1_1 = n97_O_12_1_1; // @[Top.scala 148:12]
  assign n106_I_12_1_2 = n97_O_12_1_2; // @[Top.scala 148:12]
  assign n106_I_12_2_0 = n97_O_12_2_0; // @[Top.scala 148:12]
  assign n106_I_12_2_1 = n97_O_12_2_1; // @[Top.scala 148:12]
  assign n106_I_12_2_2 = n97_O_12_2_2; // @[Top.scala 148:12]
  assign n106_I_13_0_0 = n97_O_13_0_0; // @[Top.scala 148:12]
  assign n106_I_13_0_1 = n97_O_13_0_1; // @[Top.scala 148:12]
  assign n106_I_13_0_2 = n97_O_13_0_2; // @[Top.scala 148:12]
  assign n106_I_13_1_0 = n97_O_13_1_0; // @[Top.scala 148:12]
  assign n106_I_13_1_1 = n97_O_13_1_1; // @[Top.scala 148:12]
  assign n106_I_13_1_2 = n97_O_13_1_2; // @[Top.scala 148:12]
  assign n106_I_13_2_0 = n97_O_13_2_0; // @[Top.scala 148:12]
  assign n106_I_13_2_1 = n97_O_13_2_1; // @[Top.scala 148:12]
  assign n106_I_13_2_2 = n97_O_13_2_2; // @[Top.scala 148:12]
  assign n106_I_14_0_0 = n97_O_14_0_0; // @[Top.scala 148:12]
  assign n106_I_14_0_1 = n97_O_14_0_1; // @[Top.scala 148:12]
  assign n106_I_14_0_2 = n97_O_14_0_2; // @[Top.scala 148:12]
  assign n106_I_14_1_0 = n97_O_14_1_0; // @[Top.scala 148:12]
  assign n106_I_14_1_1 = n97_O_14_1_1; // @[Top.scala 148:12]
  assign n106_I_14_1_2 = n97_O_14_1_2; // @[Top.scala 148:12]
  assign n106_I_14_2_0 = n97_O_14_2_0; // @[Top.scala 148:12]
  assign n106_I_14_2_1 = n97_O_14_2_1; // @[Top.scala 148:12]
  assign n106_I_14_2_2 = n97_O_14_2_2; // @[Top.scala 148:12]
  assign n106_I_15_0_0 = n97_O_15_0_0; // @[Top.scala 148:12]
  assign n106_I_15_0_1 = n97_O_15_0_1; // @[Top.scala 148:12]
  assign n106_I_15_0_2 = n97_O_15_0_2; // @[Top.scala 148:12]
  assign n106_I_15_1_0 = n97_O_15_1_0; // @[Top.scala 148:12]
  assign n106_I_15_1_1 = n97_O_15_1_1; // @[Top.scala 148:12]
  assign n106_I_15_1_2 = n97_O_15_1_2; // @[Top.scala 148:12]
  assign n106_I_15_2_0 = n97_O_15_2_0; // @[Top.scala 148:12]
  assign n106_I_15_2_1 = n97_O_15_2_1; // @[Top.scala 148:12]
  assign n106_I_15_2_2 = n97_O_15_2_2; // @[Top.scala 148:12]
  assign n113_valid_up = n106_valid_down; // @[Top.scala 152:19]
  assign n113_I_0_0_0_0 = n106_O_0_0_0_0; // @[Top.scala 151:12]
  assign n113_I_0_0_0_1 = n106_O_0_0_0_1; // @[Top.scala 151:12]
  assign n113_I_0_0_0_2 = n106_O_0_0_0_2; // @[Top.scala 151:12]
  assign n113_I_0_0_1_0 = n106_O_0_0_1_0; // @[Top.scala 151:12]
  assign n113_I_0_0_1_1 = n106_O_0_0_1_1; // @[Top.scala 151:12]
  assign n113_I_0_0_1_2 = n106_O_0_0_1_2; // @[Top.scala 151:12]
  assign n113_I_0_0_2_0 = n106_O_0_0_2_0; // @[Top.scala 151:12]
  assign n113_I_0_0_2_1 = n106_O_0_0_2_1; // @[Top.scala 151:12]
  assign n113_I_0_0_2_2 = n106_O_0_0_2_2; // @[Top.scala 151:12]
  assign n113_I_1_0_0_0 = n106_O_1_0_0_0; // @[Top.scala 151:12]
  assign n113_I_1_0_0_1 = n106_O_1_0_0_1; // @[Top.scala 151:12]
  assign n113_I_1_0_0_2 = n106_O_1_0_0_2; // @[Top.scala 151:12]
  assign n113_I_1_0_1_0 = n106_O_1_0_1_0; // @[Top.scala 151:12]
  assign n113_I_1_0_1_1 = n106_O_1_0_1_1; // @[Top.scala 151:12]
  assign n113_I_1_0_1_2 = n106_O_1_0_1_2; // @[Top.scala 151:12]
  assign n113_I_1_0_2_0 = n106_O_1_0_2_0; // @[Top.scala 151:12]
  assign n113_I_1_0_2_1 = n106_O_1_0_2_1; // @[Top.scala 151:12]
  assign n113_I_1_0_2_2 = n106_O_1_0_2_2; // @[Top.scala 151:12]
  assign n113_I_2_0_0_0 = n106_O_2_0_0_0; // @[Top.scala 151:12]
  assign n113_I_2_0_0_1 = n106_O_2_0_0_1; // @[Top.scala 151:12]
  assign n113_I_2_0_0_2 = n106_O_2_0_0_2; // @[Top.scala 151:12]
  assign n113_I_2_0_1_0 = n106_O_2_0_1_0; // @[Top.scala 151:12]
  assign n113_I_2_0_1_1 = n106_O_2_0_1_1; // @[Top.scala 151:12]
  assign n113_I_2_0_1_2 = n106_O_2_0_1_2; // @[Top.scala 151:12]
  assign n113_I_2_0_2_0 = n106_O_2_0_2_0; // @[Top.scala 151:12]
  assign n113_I_2_0_2_1 = n106_O_2_0_2_1; // @[Top.scala 151:12]
  assign n113_I_2_0_2_2 = n106_O_2_0_2_2; // @[Top.scala 151:12]
  assign n113_I_3_0_0_0 = n106_O_3_0_0_0; // @[Top.scala 151:12]
  assign n113_I_3_0_0_1 = n106_O_3_0_0_1; // @[Top.scala 151:12]
  assign n113_I_3_0_0_2 = n106_O_3_0_0_2; // @[Top.scala 151:12]
  assign n113_I_3_0_1_0 = n106_O_3_0_1_0; // @[Top.scala 151:12]
  assign n113_I_3_0_1_1 = n106_O_3_0_1_1; // @[Top.scala 151:12]
  assign n113_I_3_0_1_2 = n106_O_3_0_1_2; // @[Top.scala 151:12]
  assign n113_I_3_0_2_0 = n106_O_3_0_2_0; // @[Top.scala 151:12]
  assign n113_I_3_0_2_1 = n106_O_3_0_2_1; // @[Top.scala 151:12]
  assign n113_I_3_0_2_2 = n106_O_3_0_2_2; // @[Top.scala 151:12]
  assign n113_I_4_0_0_0 = n106_O_4_0_0_0; // @[Top.scala 151:12]
  assign n113_I_4_0_0_1 = n106_O_4_0_0_1; // @[Top.scala 151:12]
  assign n113_I_4_0_0_2 = n106_O_4_0_0_2; // @[Top.scala 151:12]
  assign n113_I_4_0_1_0 = n106_O_4_0_1_0; // @[Top.scala 151:12]
  assign n113_I_4_0_1_1 = n106_O_4_0_1_1; // @[Top.scala 151:12]
  assign n113_I_4_0_1_2 = n106_O_4_0_1_2; // @[Top.scala 151:12]
  assign n113_I_4_0_2_0 = n106_O_4_0_2_0; // @[Top.scala 151:12]
  assign n113_I_4_0_2_1 = n106_O_4_0_2_1; // @[Top.scala 151:12]
  assign n113_I_4_0_2_2 = n106_O_4_0_2_2; // @[Top.scala 151:12]
  assign n113_I_5_0_0_0 = n106_O_5_0_0_0; // @[Top.scala 151:12]
  assign n113_I_5_0_0_1 = n106_O_5_0_0_1; // @[Top.scala 151:12]
  assign n113_I_5_0_0_2 = n106_O_5_0_0_2; // @[Top.scala 151:12]
  assign n113_I_5_0_1_0 = n106_O_5_0_1_0; // @[Top.scala 151:12]
  assign n113_I_5_0_1_1 = n106_O_5_0_1_1; // @[Top.scala 151:12]
  assign n113_I_5_0_1_2 = n106_O_5_0_1_2; // @[Top.scala 151:12]
  assign n113_I_5_0_2_0 = n106_O_5_0_2_0; // @[Top.scala 151:12]
  assign n113_I_5_0_2_1 = n106_O_5_0_2_1; // @[Top.scala 151:12]
  assign n113_I_5_0_2_2 = n106_O_5_0_2_2; // @[Top.scala 151:12]
  assign n113_I_6_0_0_0 = n106_O_6_0_0_0; // @[Top.scala 151:12]
  assign n113_I_6_0_0_1 = n106_O_6_0_0_1; // @[Top.scala 151:12]
  assign n113_I_6_0_0_2 = n106_O_6_0_0_2; // @[Top.scala 151:12]
  assign n113_I_6_0_1_0 = n106_O_6_0_1_0; // @[Top.scala 151:12]
  assign n113_I_6_0_1_1 = n106_O_6_0_1_1; // @[Top.scala 151:12]
  assign n113_I_6_0_1_2 = n106_O_6_0_1_2; // @[Top.scala 151:12]
  assign n113_I_6_0_2_0 = n106_O_6_0_2_0; // @[Top.scala 151:12]
  assign n113_I_6_0_2_1 = n106_O_6_0_2_1; // @[Top.scala 151:12]
  assign n113_I_6_0_2_2 = n106_O_6_0_2_2; // @[Top.scala 151:12]
  assign n113_I_7_0_0_0 = n106_O_7_0_0_0; // @[Top.scala 151:12]
  assign n113_I_7_0_0_1 = n106_O_7_0_0_1; // @[Top.scala 151:12]
  assign n113_I_7_0_0_2 = n106_O_7_0_0_2; // @[Top.scala 151:12]
  assign n113_I_7_0_1_0 = n106_O_7_0_1_0; // @[Top.scala 151:12]
  assign n113_I_7_0_1_1 = n106_O_7_0_1_1; // @[Top.scala 151:12]
  assign n113_I_7_0_1_2 = n106_O_7_0_1_2; // @[Top.scala 151:12]
  assign n113_I_7_0_2_0 = n106_O_7_0_2_0; // @[Top.scala 151:12]
  assign n113_I_7_0_2_1 = n106_O_7_0_2_1; // @[Top.scala 151:12]
  assign n113_I_7_0_2_2 = n106_O_7_0_2_2; // @[Top.scala 151:12]
  assign n113_I_8_0_0_0 = n106_O_8_0_0_0; // @[Top.scala 151:12]
  assign n113_I_8_0_0_1 = n106_O_8_0_0_1; // @[Top.scala 151:12]
  assign n113_I_8_0_0_2 = n106_O_8_0_0_2; // @[Top.scala 151:12]
  assign n113_I_8_0_1_0 = n106_O_8_0_1_0; // @[Top.scala 151:12]
  assign n113_I_8_0_1_1 = n106_O_8_0_1_1; // @[Top.scala 151:12]
  assign n113_I_8_0_1_2 = n106_O_8_0_1_2; // @[Top.scala 151:12]
  assign n113_I_8_0_2_0 = n106_O_8_0_2_0; // @[Top.scala 151:12]
  assign n113_I_8_0_2_1 = n106_O_8_0_2_1; // @[Top.scala 151:12]
  assign n113_I_8_0_2_2 = n106_O_8_0_2_2; // @[Top.scala 151:12]
  assign n113_I_9_0_0_0 = n106_O_9_0_0_0; // @[Top.scala 151:12]
  assign n113_I_9_0_0_1 = n106_O_9_0_0_1; // @[Top.scala 151:12]
  assign n113_I_9_0_0_2 = n106_O_9_0_0_2; // @[Top.scala 151:12]
  assign n113_I_9_0_1_0 = n106_O_9_0_1_0; // @[Top.scala 151:12]
  assign n113_I_9_0_1_1 = n106_O_9_0_1_1; // @[Top.scala 151:12]
  assign n113_I_9_0_1_2 = n106_O_9_0_1_2; // @[Top.scala 151:12]
  assign n113_I_9_0_2_0 = n106_O_9_0_2_0; // @[Top.scala 151:12]
  assign n113_I_9_0_2_1 = n106_O_9_0_2_1; // @[Top.scala 151:12]
  assign n113_I_9_0_2_2 = n106_O_9_0_2_2; // @[Top.scala 151:12]
  assign n113_I_10_0_0_0 = n106_O_10_0_0_0; // @[Top.scala 151:12]
  assign n113_I_10_0_0_1 = n106_O_10_0_0_1; // @[Top.scala 151:12]
  assign n113_I_10_0_0_2 = n106_O_10_0_0_2; // @[Top.scala 151:12]
  assign n113_I_10_0_1_0 = n106_O_10_0_1_0; // @[Top.scala 151:12]
  assign n113_I_10_0_1_1 = n106_O_10_0_1_1; // @[Top.scala 151:12]
  assign n113_I_10_0_1_2 = n106_O_10_0_1_2; // @[Top.scala 151:12]
  assign n113_I_10_0_2_0 = n106_O_10_0_2_0; // @[Top.scala 151:12]
  assign n113_I_10_0_2_1 = n106_O_10_0_2_1; // @[Top.scala 151:12]
  assign n113_I_10_0_2_2 = n106_O_10_0_2_2; // @[Top.scala 151:12]
  assign n113_I_11_0_0_0 = n106_O_11_0_0_0; // @[Top.scala 151:12]
  assign n113_I_11_0_0_1 = n106_O_11_0_0_1; // @[Top.scala 151:12]
  assign n113_I_11_0_0_2 = n106_O_11_0_0_2; // @[Top.scala 151:12]
  assign n113_I_11_0_1_0 = n106_O_11_0_1_0; // @[Top.scala 151:12]
  assign n113_I_11_0_1_1 = n106_O_11_0_1_1; // @[Top.scala 151:12]
  assign n113_I_11_0_1_2 = n106_O_11_0_1_2; // @[Top.scala 151:12]
  assign n113_I_11_0_2_0 = n106_O_11_0_2_0; // @[Top.scala 151:12]
  assign n113_I_11_0_2_1 = n106_O_11_0_2_1; // @[Top.scala 151:12]
  assign n113_I_11_0_2_2 = n106_O_11_0_2_2; // @[Top.scala 151:12]
  assign n113_I_12_0_0_0 = n106_O_12_0_0_0; // @[Top.scala 151:12]
  assign n113_I_12_0_0_1 = n106_O_12_0_0_1; // @[Top.scala 151:12]
  assign n113_I_12_0_0_2 = n106_O_12_0_0_2; // @[Top.scala 151:12]
  assign n113_I_12_0_1_0 = n106_O_12_0_1_0; // @[Top.scala 151:12]
  assign n113_I_12_0_1_1 = n106_O_12_0_1_1; // @[Top.scala 151:12]
  assign n113_I_12_0_1_2 = n106_O_12_0_1_2; // @[Top.scala 151:12]
  assign n113_I_12_0_2_0 = n106_O_12_0_2_0; // @[Top.scala 151:12]
  assign n113_I_12_0_2_1 = n106_O_12_0_2_1; // @[Top.scala 151:12]
  assign n113_I_12_0_2_2 = n106_O_12_0_2_2; // @[Top.scala 151:12]
  assign n113_I_13_0_0_0 = n106_O_13_0_0_0; // @[Top.scala 151:12]
  assign n113_I_13_0_0_1 = n106_O_13_0_0_1; // @[Top.scala 151:12]
  assign n113_I_13_0_0_2 = n106_O_13_0_0_2; // @[Top.scala 151:12]
  assign n113_I_13_0_1_0 = n106_O_13_0_1_0; // @[Top.scala 151:12]
  assign n113_I_13_0_1_1 = n106_O_13_0_1_1; // @[Top.scala 151:12]
  assign n113_I_13_0_1_2 = n106_O_13_0_1_2; // @[Top.scala 151:12]
  assign n113_I_13_0_2_0 = n106_O_13_0_2_0; // @[Top.scala 151:12]
  assign n113_I_13_0_2_1 = n106_O_13_0_2_1; // @[Top.scala 151:12]
  assign n113_I_13_0_2_2 = n106_O_13_0_2_2; // @[Top.scala 151:12]
  assign n113_I_14_0_0_0 = n106_O_14_0_0_0; // @[Top.scala 151:12]
  assign n113_I_14_0_0_1 = n106_O_14_0_0_1; // @[Top.scala 151:12]
  assign n113_I_14_0_0_2 = n106_O_14_0_0_2; // @[Top.scala 151:12]
  assign n113_I_14_0_1_0 = n106_O_14_0_1_0; // @[Top.scala 151:12]
  assign n113_I_14_0_1_1 = n106_O_14_0_1_1; // @[Top.scala 151:12]
  assign n113_I_14_0_1_2 = n106_O_14_0_1_2; // @[Top.scala 151:12]
  assign n113_I_14_0_2_0 = n106_O_14_0_2_0; // @[Top.scala 151:12]
  assign n113_I_14_0_2_1 = n106_O_14_0_2_1; // @[Top.scala 151:12]
  assign n113_I_14_0_2_2 = n106_O_14_0_2_2; // @[Top.scala 151:12]
  assign n113_I_15_0_0_0 = n106_O_15_0_0_0; // @[Top.scala 151:12]
  assign n113_I_15_0_0_1 = n106_O_15_0_0_1; // @[Top.scala 151:12]
  assign n113_I_15_0_0_2 = n106_O_15_0_0_2; // @[Top.scala 151:12]
  assign n113_I_15_0_1_0 = n106_O_15_0_1_0; // @[Top.scala 151:12]
  assign n113_I_15_0_1_1 = n106_O_15_0_1_1; // @[Top.scala 151:12]
  assign n113_I_15_0_1_2 = n106_O_15_0_1_2; // @[Top.scala 151:12]
  assign n113_I_15_0_2_0 = n106_O_15_0_2_0; // @[Top.scala 151:12]
  assign n113_I_15_0_2_1 = n106_O_15_0_2_1; // @[Top.scala 151:12]
  assign n113_I_15_0_2_2 = n106_O_15_0_2_2; // @[Top.scala 151:12]
  assign n155_clock = clock;
  assign n155_reset = reset;
  assign n155_valid_up = n113_valid_down; // @[Top.scala 155:19]
  assign n155_I_0_0_0 = n113_O_0_0_0; // @[Top.scala 154:12]
  assign n155_I_0_0_1 = n113_O_0_0_1; // @[Top.scala 154:12]
  assign n155_I_0_0_2 = n113_O_0_0_2; // @[Top.scala 154:12]
  assign n155_I_0_1_0 = n113_O_0_1_0; // @[Top.scala 154:12]
  assign n155_I_0_1_1 = n113_O_0_1_1; // @[Top.scala 154:12]
  assign n155_I_0_1_2 = n113_O_0_1_2; // @[Top.scala 154:12]
  assign n155_I_0_2_0 = n113_O_0_2_0; // @[Top.scala 154:12]
  assign n155_I_0_2_1 = n113_O_0_2_1; // @[Top.scala 154:12]
  assign n155_I_0_2_2 = n113_O_0_2_2; // @[Top.scala 154:12]
  assign n155_I_1_0_0 = n113_O_1_0_0; // @[Top.scala 154:12]
  assign n155_I_1_0_1 = n113_O_1_0_1; // @[Top.scala 154:12]
  assign n155_I_1_0_2 = n113_O_1_0_2; // @[Top.scala 154:12]
  assign n155_I_1_1_0 = n113_O_1_1_0; // @[Top.scala 154:12]
  assign n155_I_1_1_1 = n113_O_1_1_1; // @[Top.scala 154:12]
  assign n155_I_1_1_2 = n113_O_1_1_2; // @[Top.scala 154:12]
  assign n155_I_1_2_0 = n113_O_1_2_0; // @[Top.scala 154:12]
  assign n155_I_1_2_1 = n113_O_1_2_1; // @[Top.scala 154:12]
  assign n155_I_1_2_2 = n113_O_1_2_2; // @[Top.scala 154:12]
  assign n155_I_2_0_0 = n113_O_2_0_0; // @[Top.scala 154:12]
  assign n155_I_2_0_1 = n113_O_2_0_1; // @[Top.scala 154:12]
  assign n155_I_2_0_2 = n113_O_2_0_2; // @[Top.scala 154:12]
  assign n155_I_2_1_0 = n113_O_2_1_0; // @[Top.scala 154:12]
  assign n155_I_2_1_1 = n113_O_2_1_1; // @[Top.scala 154:12]
  assign n155_I_2_1_2 = n113_O_2_1_2; // @[Top.scala 154:12]
  assign n155_I_2_2_0 = n113_O_2_2_0; // @[Top.scala 154:12]
  assign n155_I_2_2_1 = n113_O_2_2_1; // @[Top.scala 154:12]
  assign n155_I_2_2_2 = n113_O_2_2_2; // @[Top.scala 154:12]
  assign n155_I_3_0_0 = n113_O_3_0_0; // @[Top.scala 154:12]
  assign n155_I_3_0_1 = n113_O_3_0_1; // @[Top.scala 154:12]
  assign n155_I_3_0_2 = n113_O_3_0_2; // @[Top.scala 154:12]
  assign n155_I_3_1_0 = n113_O_3_1_0; // @[Top.scala 154:12]
  assign n155_I_3_1_1 = n113_O_3_1_1; // @[Top.scala 154:12]
  assign n155_I_3_1_2 = n113_O_3_1_2; // @[Top.scala 154:12]
  assign n155_I_3_2_0 = n113_O_3_2_0; // @[Top.scala 154:12]
  assign n155_I_3_2_1 = n113_O_3_2_1; // @[Top.scala 154:12]
  assign n155_I_3_2_2 = n113_O_3_2_2; // @[Top.scala 154:12]
  assign n155_I_4_0_0 = n113_O_4_0_0; // @[Top.scala 154:12]
  assign n155_I_4_0_1 = n113_O_4_0_1; // @[Top.scala 154:12]
  assign n155_I_4_0_2 = n113_O_4_0_2; // @[Top.scala 154:12]
  assign n155_I_4_1_0 = n113_O_4_1_0; // @[Top.scala 154:12]
  assign n155_I_4_1_1 = n113_O_4_1_1; // @[Top.scala 154:12]
  assign n155_I_4_1_2 = n113_O_4_1_2; // @[Top.scala 154:12]
  assign n155_I_4_2_0 = n113_O_4_2_0; // @[Top.scala 154:12]
  assign n155_I_4_2_1 = n113_O_4_2_1; // @[Top.scala 154:12]
  assign n155_I_4_2_2 = n113_O_4_2_2; // @[Top.scala 154:12]
  assign n155_I_5_0_0 = n113_O_5_0_0; // @[Top.scala 154:12]
  assign n155_I_5_0_1 = n113_O_5_0_1; // @[Top.scala 154:12]
  assign n155_I_5_0_2 = n113_O_5_0_2; // @[Top.scala 154:12]
  assign n155_I_5_1_0 = n113_O_5_1_0; // @[Top.scala 154:12]
  assign n155_I_5_1_1 = n113_O_5_1_1; // @[Top.scala 154:12]
  assign n155_I_5_1_2 = n113_O_5_1_2; // @[Top.scala 154:12]
  assign n155_I_5_2_0 = n113_O_5_2_0; // @[Top.scala 154:12]
  assign n155_I_5_2_1 = n113_O_5_2_1; // @[Top.scala 154:12]
  assign n155_I_5_2_2 = n113_O_5_2_2; // @[Top.scala 154:12]
  assign n155_I_6_0_0 = n113_O_6_0_0; // @[Top.scala 154:12]
  assign n155_I_6_0_1 = n113_O_6_0_1; // @[Top.scala 154:12]
  assign n155_I_6_0_2 = n113_O_6_0_2; // @[Top.scala 154:12]
  assign n155_I_6_1_0 = n113_O_6_1_0; // @[Top.scala 154:12]
  assign n155_I_6_1_1 = n113_O_6_1_1; // @[Top.scala 154:12]
  assign n155_I_6_1_2 = n113_O_6_1_2; // @[Top.scala 154:12]
  assign n155_I_6_2_0 = n113_O_6_2_0; // @[Top.scala 154:12]
  assign n155_I_6_2_1 = n113_O_6_2_1; // @[Top.scala 154:12]
  assign n155_I_6_2_2 = n113_O_6_2_2; // @[Top.scala 154:12]
  assign n155_I_7_0_0 = n113_O_7_0_0; // @[Top.scala 154:12]
  assign n155_I_7_0_1 = n113_O_7_0_1; // @[Top.scala 154:12]
  assign n155_I_7_0_2 = n113_O_7_0_2; // @[Top.scala 154:12]
  assign n155_I_7_1_0 = n113_O_7_1_0; // @[Top.scala 154:12]
  assign n155_I_7_1_1 = n113_O_7_1_1; // @[Top.scala 154:12]
  assign n155_I_7_1_2 = n113_O_7_1_2; // @[Top.scala 154:12]
  assign n155_I_7_2_0 = n113_O_7_2_0; // @[Top.scala 154:12]
  assign n155_I_7_2_1 = n113_O_7_2_1; // @[Top.scala 154:12]
  assign n155_I_7_2_2 = n113_O_7_2_2; // @[Top.scala 154:12]
  assign n155_I_8_0_0 = n113_O_8_0_0; // @[Top.scala 154:12]
  assign n155_I_8_0_1 = n113_O_8_0_1; // @[Top.scala 154:12]
  assign n155_I_8_0_2 = n113_O_8_0_2; // @[Top.scala 154:12]
  assign n155_I_8_1_0 = n113_O_8_1_0; // @[Top.scala 154:12]
  assign n155_I_8_1_1 = n113_O_8_1_1; // @[Top.scala 154:12]
  assign n155_I_8_1_2 = n113_O_8_1_2; // @[Top.scala 154:12]
  assign n155_I_8_2_0 = n113_O_8_2_0; // @[Top.scala 154:12]
  assign n155_I_8_2_1 = n113_O_8_2_1; // @[Top.scala 154:12]
  assign n155_I_8_2_2 = n113_O_8_2_2; // @[Top.scala 154:12]
  assign n155_I_9_0_0 = n113_O_9_0_0; // @[Top.scala 154:12]
  assign n155_I_9_0_1 = n113_O_9_0_1; // @[Top.scala 154:12]
  assign n155_I_9_0_2 = n113_O_9_0_2; // @[Top.scala 154:12]
  assign n155_I_9_1_0 = n113_O_9_1_0; // @[Top.scala 154:12]
  assign n155_I_9_1_1 = n113_O_9_1_1; // @[Top.scala 154:12]
  assign n155_I_9_1_2 = n113_O_9_1_2; // @[Top.scala 154:12]
  assign n155_I_9_2_0 = n113_O_9_2_0; // @[Top.scala 154:12]
  assign n155_I_9_2_1 = n113_O_9_2_1; // @[Top.scala 154:12]
  assign n155_I_9_2_2 = n113_O_9_2_2; // @[Top.scala 154:12]
  assign n155_I_10_0_0 = n113_O_10_0_0; // @[Top.scala 154:12]
  assign n155_I_10_0_1 = n113_O_10_0_1; // @[Top.scala 154:12]
  assign n155_I_10_0_2 = n113_O_10_0_2; // @[Top.scala 154:12]
  assign n155_I_10_1_0 = n113_O_10_1_0; // @[Top.scala 154:12]
  assign n155_I_10_1_1 = n113_O_10_1_1; // @[Top.scala 154:12]
  assign n155_I_10_1_2 = n113_O_10_1_2; // @[Top.scala 154:12]
  assign n155_I_10_2_0 = n113_O_10_2_0; // @[Top.scala 154:12]
  assign n155_I_10_2_1 = n113_O_10_2_1; // @[Top.scala 154:12]
  assign n155_I_10_2_2 = n113_O_10_2_2; // @[Top.scala 154:12]
  assign n155_I_11_0_0 = n113_O_11_0_0; // @[Top.scala 154:12]
  assign n155_I_11_0_1 = n113_O_11_0_1; // @[Top.scala 154:12]
  assign n155_I_11_0_2 = n113_O_11_0_2; // @[Top.scala 154:12]
  assign n155_I_11_1_0 = n113_O_11_1_0; // @[Top.scala 154:12]
  assign n155_I_11_1_1 = n113_O_11_1_1; // @[Top.scala 154:12]
  assign n155_I_11_1_2 = n113_O_11_1_2; // @[Top.scala 154:12]
  assign n155_I_11_2_0 = n113_O_11_2_0; // @[Top.scala 154:12]
  assign n155_I_11_2_1 = n113_O_11_2_1; // @[Top.scala 154:12]
  assign n155_I_11_2_2 = n113_O_11_2_2; // @[Top.scala 154:12]
  assign n155_I_12_0_0 = n113_O_12_0_0; // @[Top.scala 154:12]
  assign n155_I_12_0_1 = n113_O_12_0_1; // @[Top.scala 154:12]
  assign n155_I_12_0_2 = n113_O_12_0_2; // @[Top.scala 154:12]
  assign n155_I_12_1_0 = n113_O_12_1_0; // @[Top.scala 154:12]
  assign n155_I_12_1_1 = n113_O_12_1_1; // @[Top.scala 154:12]
  assign n155_I_12_1_2 = n113_O_12_1_2; // @[Top.scala 154:12]
  assign n155_I_12_2_0 = n113_O_12_2_0; // @[Top.scala 154:12]
  assign n155_I_12_2_1 = n113_O_12_2_1; // @[Top.scala 154:12]
  assign n155_I_12_2_2 = n113_O_12_2_2; // @[Top.scala 154:12]
  assign n155_I_13_0_0 = n113_O_13_0_0; // @[Top.scala 154:12]
  assign n155_I_13_0_1 = n113_O_13_0_1; // @[Top.scala 154:12]
  assign n155_I_13_0_2 = n113_O_13_0_2; // @[Top.scala 154:12]
  assign n155_I_13_1_0 = n113_O_13_1_0; // @[Top.scala 154:12]
  assign n155_I_13_1_1 = n113_O_13_1_1; // @[Top.scala 154:12]
  assign n155_I_13_1_2 = n113_O_13_1_2; // @[Top.scala 154:12]
  assign n155_I_13_2_0 = n113_O_13_2_0; // @[Top.scala 154:12]
  assign n155_I_13_2_1 = n113_O_13_2_1; // @[Top.scala 154:12]
  assign n155_I_13_2_2 = n113_O_13_2_2; // @[Top.scala 154:12]
  assign n155_I_14_0_0 = n113_O_14_0_0; // @[Top.scala 154:12]
  assign n155_I_14_0_1 = n113_O_14_0_1; // @[Top.scala 154:12]
  assign n155_I_14_0_2 = n113_O_14_0_2; // @[Top.scala 154:12]
  assign n155_I_14_1_0 = n113_O_14_1_0; // @[Top.scala 154:12]
  assign n155_I_14_1_1 = n113_O_14_1_1; // @[Top.scala 154:12]
  assign n155_I_14_1_2 = n113_O_14_1_2; // @[Top.scala 154:12]
  assign n155_I_14_2_0 = n113_O_14_2_0; // @[Top.scala 154:12]
  assign n155_I_14_2_1 = n113_O_14_2_1; // @[Top.scala 154:12]
  assign n155_I_14_2_2 = n113_O_14_2_2; // @[Top.scala 154:12]
  assign n155_I_15_0_0 = n113_O_15_0_0; // @[Top.scala 154:12]
  assign n155_I_15_0_1 = n113_O_15_0_1; // @[Top.scala 154:12]
  assign n155_I_15_0_2 = n113_O_15_0_2; // @[Top.scala 154:12]
  assign n155_I_15_1_0 = n113_O_15_1_0; // @[Top.scala 154:12]
  assign n155_I_15_1_1 = n113_O_15_1_1; // @[Top.scala 154:12]
  assign n155_I_15_1_2 = n113_O_15_1_2; // @[Top.scala 154:12]
  assign n155_I_15_2_0 = n113_O_15_2_0; // @[Top.scala 154:12]
  assign n155_I_15_2_1 = n113_O_15_2_1; // @[Top.scala 154:12]
  assign n155_I_15_2_2 = n113_O_15_2_2; // @[Top.scala 154:12]
  assign n156_valid_up = n155_valid_down; // @[Top.scala 158:19]
  assign n156_I_0_0_0 = n155_O_0_0_0; // @[Top.scala 157:12]
  assign n156_I_1_0_0 = n155_O_1_0_0; // @[Top.scala 157:12]
  assign n156_I_2_0_0 = n155_O_2_0_0; // @[Top.scala 157:12]
  assign n156_I_3_0_0 = n155_O_3_0_0; // @[Top.scala 157:12]
  assign n156_I_4_0_0 = n155_O_4_0_0; // @[Top.scala 157:12]
  assign n156_I_5_0_0 = n155_O_5_0_0; // @[Top.scala 157:12]
  assign n156_I_6_0_0 = n155_O_6_0_0; // @[Top.scala 157:12]
  assign n156_I_7_0_0 = n155_O_7_0_0; // @[Top.scala 157:12]
  assign n156_I_8_0_0 = n155_O_8_0_0; // @[Top.scala 157:12]
  assign n156_I_9_0_0 = n155_O_9_0_0; // @[Top.scala 157:12]
  assign n156_I_10_0_0 = n155_O_10_0_0; // @[Top.scala 157:12]
  assign n156_I_11_0_0 = n155_O_11_0_0; // @[Top.scala 157:12]
  assign n156_I_12_0_0 = n155_O_12_0_0; // @[Top.scala 157:12]
  assign n156_I_13_0_0 = n155_O_13_0_0; // @[Top.scala 157:12]
  assign n156_I_14_0_0 = n155_O_14_0_0; // @[Top.scala 157:12]
  assign n156_I_15_0_0 = n155_O_15_0_0; // @[Top.scala 157:12]
  assign n157_valid_up = n156_valid_down; // @[Top.scala 161:19]
  assign n157_I_0_0 = n156_O_0_0; // @[Top.scala 160:12]
  assign n157_I_1_0 = n156_O_1_0; // @[Top.scala 160:12]
  assign n157_I_2_0 = n156_O_2_0; // @[Top.scala 160:12]
  assign n157_I_3_0 = n156_O_3_0; // @[Top.scala 160:12]
  assign n157_I_4_0 = n156_O_4_0; // @[Top.scala 160:12]
  assign n157_I_5_0 = n156_O_5_0; // @[Top.scala 160:12]
  assign n157_I_6_0 = n156_O_6_0; // @[Top.scala 160:12]
  assign n157_I_7_0 = n156_O_7_0; // @[Top.scala 160:12]
  assign n157_I_8_0 = n156_O_8_0; // @[Top.scala 160:12]
  assign n157_I_9_0 = n156_O_9_0; // @[Top.scala 160:12]
  assign n157_I_10_0 = n156_O_10_0; // @[Top.scala 160:12]
  assign n157_I_11_0 = n156_O_11_0; // @[Top.scala 160:12]
  assign n157_I_12_0 = n156_O_12_0; // @[Top.scala 160:12]
  assign n157_I_13_0 = n156_O_13_0; // @[Top.scala 160:12]
  assign n157_I_14_0 = n156_O_14_0; // @[Top.scala 160:12]
  assign n157_I_15_0 = n156_O_15_0; // @[Top.scala 160:12]
  assign n158_clock = clock;
  assign n158_reset = reset;
  assign n158_valid_up = n157_valid_down; // @[Top.scala 164:19]
  assign n158_I_0 = n157_O_0; // @[Top.scala 163:12]
  assign n158_I_1 = n157_O_1; // @[Top.scala 163:12]
  assign n158_I_2 = n157_O_2; // @[Top.scala 163:12]
  assign n158_I_3 = n157_O_3; // @[Top.scala 163:12]
  assign n158_I_4 = n157_O_4; // @[Top.scala 163:12]
  assign n158_I_5 = n157_O_5; // @[Top.scala 163:12]
  assign n158_I_6 = n157_O_6; // @[Top.scala 163:12]
  assign n158_I_7 = n157_O_7; // @[Top.scala 163:12]
  assign n158_I_8 = n157_O_8; // @[Top.scala 163:12]
  assign n158_I_9 = n157_O_9; // @[Top.scala 163:12]
  assign n158_I_10 = n157_O_10; // @[Top.scala 163:12]
  assign n158_I_11 = n157_O_11; // @[Top.scala 163:12]
  assign n158_I_12 = n157_O_12; // @[Top.scala 163:12]
  assign n158_I_13 = n157_O_13; // @[Top.scala 163:12]
  assign n158_I_14 = n157_O_14; // @[Top.scala 163:12]
  assign n158_I_15 = n157_O_15; // @[Top.scala 163:12]
  assign n159_clock = clock;
  assign n159_reset = reset;
  assign n159_valid_up = n158_valid_down; // @[Top.scala 167:19]
  assign n159_I_0 = n158_O_0; // @[Top.scala 166:12]
  assign n159_I_1 = n158_O_1; // @[Top.scala 166:12]
  assign n159_I_2 = n158_O_2; // @[Top.scala 166:12]
  assign n159_I_3 = n158_O_3; // @[Top.scala 166:12]
  assign n159_I_4 = n158_O_4; // @[Top.scala 166:12]
  assign n159_I_5 = n158_O_5; // @[Top.scala 166:12]
  assign n159_I_6 = n158_O_6; // @[Top.scala 166:12]
  assign n159_I_7 = n158_O_7; // @[Top.scala 166:12]
  assign n159_I_8 = n158_O_8; // @[Top.scala 166:12]
  assign n159_I_9 = n158_O_9; // @[Top.scala 166:12]
  assign n159_I_10 = n158_O_10; // @[Top.scala 166:12]
  assign n159_I_11 = n158_O_11; // @[Top.scala 166:12]
  assign n159_I_12 = n158_O_12; // @[Top.scala 166:12]
  assign n159_I_13 = n158_O_13; // @[Top.scala 166:12]
  assign n159_I_14 = n158_O_14; // @[Top.scala 166:12]
  assign n159_I_15 = n158_O_15; // @[Top.scala 166:12]
  assign n160_clock = clock;
  assign n160_reset = reset;
  assign n160_valid_up = n159_valid_down; // @[Top.scala 170:19]
  assign n160_I_0 = n159_O_0; // @[Top.scala 169:12]
  assign n160_I_1 = n159_O_1; // @[Top.scala 169:12]
  assign n160_I_2 = n159_O_2; // @[Top.scala 169:12]
  assign n160_I_3 = n159_O_3; // @[Top.scala 169:12]
  assign n160_I_4 = n159_O_4; // @[Top.scala 169:12]
  assign n160_I_5 = n159_O_5; // @[Top.scala 169:12]
  assign n160_I_6 = n159_O_6; // @[Top.scala 169:12]
  assign n160_I_7 = n159_O_7; // @[Top.scala 169:12]
  assign n160_I_8 = n159_O_8; // @[Top.scala 169:12]
  assign n160_I_9 = n159_O_9; // @[Top.scala 169:12]
  assign n160_I_10 = n159_O_10; // @[Top.scala 169:12]
  assign n160_I_11 = n159_O_11; // @[Top.scala 169:12]
  assign n160_I_12 = n159_O_12; // @[Top.scala 169:12]
  assign n160_I_13 = n159_O_13; // @[Top.scala 169:12]
  assign n160_I_14 = n159_O_14; // @[Top.scala 169:12]
  assign n160_I_15 = n159_O_15; // @[Top.scala 169:12]
endmodule
