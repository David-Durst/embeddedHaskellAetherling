p// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  output [31:0] O_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x349_inr_Foreach_SAMPLER_BOX_kernelx349_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x194_TREADY(dontcare), // @[:@1298.4]
    .io_in_x194_TDATA(I_0), // @[:@1298.4]
    .io_in_x194_TID(8'h0),
    .io_in_x194_TDEST(8'h0),
    .io_in_x195_TVALID(valid_down), // @[:@1298.4]
    .io_in_x195_TDATA(O_0), // @[:@1298.4]
    .io_in_x195_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x202_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule


// End boilerplate
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4b); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh4b); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x196_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x475_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x341_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x197_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x198_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x202_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x216_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x390_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x208_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x216_inr_Foreach_kernelx216_inr_Foreach_concrete1( // @[:@4712.2]
  input         clock, // @[:@4713.4]
  input         reset, // @[:@4714.4]
  output        io_in_x198_fifoinpacked_0_wPort_0_en_0, // @[:@4715.4]
  input         io_in_x198_fifoinpacked_0_full, // @[:@4715.4]
  output        io_in_x198_fifoinpacked_0_active_0_in, // @[:@4715.4]
  input         io_in_x198_fifoinpacked_0_active_0_out, // @[:@4715.4]
  input         io_sigsIn_backpressure, // @[:@4715.4]
  input         io_sigsIn_datapathEn, // @[:@4715.4]
  input         io_sigsIn_break, // @[:@4715.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@4715.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4715.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4715.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@4715.4]
  input         io_rr // @[:@4715.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4749.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4749.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4761.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@4761.4]
  wire  x390_sub_1_clock; // @[Math.scala 191:24:@4788.4]
  wire  x390_sub_1_reset; // @[Math.scala 191:24:@4788.4]
  wire [31:0] x390_sub_1_io_a; // @[Math.scala 191:24:@4788.4]
  wire [31:0] x390_sub_1_io_b; // @[Math.scala 191:24:@4788.4]
  wire  x390_sub_1_io_flow; // @[Math.scala 191:24:@4788.4]
  wire [31:0] x390_sub_1_io_result; // @[Math.scala 191:24:@4788.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4798.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4798.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4798.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4798.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4798.4]
  wire  x208_sum_1_clock; // @[Math.scala 150:24:@4807.4]
  wire  x208_sum_1_reset; // @[Math.scala 150:24:@4807.4]
  wire [31:0] x208_sum_1_io_a; // @[Math.scala 150:24:@4807.4]
  wire [31:0] x208_sum_1_io_b; // @[Math.scala 150:24:@4807.4]
  wire  x208_sum_1_io_flow; // @[Math.scala 150:24:@4807.4]
  wire [31:0] x208_sum_1_io_result; // @[Math.scala 150:24:@4807.4]
  wire  x209_sum_1_clock; // @[Math.scala 150:24:@4819.4]
  wire  x209_sum_1_reset; // @[Math.scala 150:24:@4819.4]
  wire [31:0] x209_sum_1_io_a; // @[Math.scala 150:24:@4819.4]
  wire [31:0] x209_sum_1_io_b; // @[Math.scala 150:24:@4819.4]
  wire  x209_sum_1_io_flow; // @[Math.scala 150:24:@4819.4]
  wire [31:0] x209_sum_1_io_result; // @[Math.scala 150:24:@4819.4]
  wire  x392_sum_1_clock; // @[Math.scala 150:24:@4834.4]
  wire  x392_sum_1_reset; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x392_sum_1_io_a; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x392_sum_1_io_b; // @[Math.scala 150:24:@4834.4]
  wire  x392_sum_1_io_flow; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x392_sum_1_io_result; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x212_1_io_b; // @[Math.scala 720:24:@4855.4]
  wire [31:0] x212_1_io_result; // @[Math.scala 720:24:@4855.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4888.4]
  wire  _T_327; // @[sm_x216_inr_Foreach.scala 62:18:@4774.4]
  wire  _T_328; // @[sm_x216_inr_Foreach.scala 62:55:@4775.4]
  wire [31:0] b203_number; // @[Math.scala 723:22:@4754.4 Math.scala 724:14:@4755.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@4779.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@4779.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@4784.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@4784.4]
  wire [31:0] x209_sum_number; // @[Math.scala 154:22:@4825.4 Math.scala 155:14:@4826.4]
  wire [33:0] _GEN_2; // @[Math.scala 461:32:@4830.4]
  wire [33:0] _T_353; // @[Math.scala 461:32:@4830.4]
  wire [31:0] x392_sum_number; // @[Math.scala 154:22:@4840.4 Math.scala 155:14:@4841.4]
  wire [31:0] _T_364; // @[Math.scala 406:49:@4847.4]
  wire [31:0] _T_366; // @[Math.scala 406:56:@4849.4]
  wire [31:0] _T_367; // @[Math.scala 406:56:@4850.4]
  wire  _T_385; // @[sm_x216_inr_Foreach.scala 93:131:@4885.4]
  wire  _T_389; // @[package.scala 96:25:@4893.4 package.scala 96:25:@4894.4]
  wire  _T_391; // @[implicits.scala 55:10:@4895.4]
  wire  _T_392; // @[sm_x216_inr_Foreach.scala 93:148:@4896.4]
  wire  _T_394; // @[sm_x216_inr_Foreach.scala 93:236:@4898.4]
  wire  _T_395; // @[sm_x216_inr_Foreach.scala 93:255:@4899.4]
  wire  x478_b205_D4; // @[package.scala 96:25:@4873.4 package.scala 96:25:@4874.4]
  wire  _T_398; // @[sm_x216_inr_Foreach.scala 93:291:@4901.4]
  wire  x479_b206_D4; // @[package.scala 96:25:@4882.4 package.scala 96:25:@4883.4]
  _ _ ( // @[Math.scala 720:24:@4749.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@4761.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x390_sub x390_sub_1 ( // @[Math.scala 191:24:@4788.4]
    .clock(x390_sub_1_clock),
    .reset(x390_sub_1_reset),
    .io_a(x390_sub_1_io_a),
    .io_b(x390_sub_1_io_b),
    .io_flow(x390_sub_1_io_flow),
    .io_result(x390_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@4798.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x208_sum x208_sum_1 ( // @[Math.scala 150:24:@4807.4]
    .clock(x208_sum_1_clock),
    .reset(x208_sum_1_reset),
    .io_a(x208_sum_1_io_a),
    .io_b(x208_sum_1_io_b),
    .io_flow(x208_sum_1_io_flow),
    .io_result(x208_sum_1_io_result)
  );
  x208_sum x209_sum_1 ( // @[Math.scala 150:24:@4819.4]
    .clock(x209_sum_1_clock),
    .reset(x209_sum_1_reset),
    .io_a(x209_sum_1_io_a),
    .io_b(x209_sum_1_io_b),
    .io_flow(x209_sum_1_io_flow),
    .io_result(x209_sum_1_io_result)
  );
  x208_sum x392_sum_1 ( // @[Math.scala 150:24:@4834.4]
    .clock(x392_sum_1_clock),
    .reset(x392_sum_1_reset),
    .io_a(x392_sum_1_io_a),
    .io_b(x392_sum_1_io_b),
    .io_flow(x392_sum_1_io_flow),
    .io_result(x392_sum_1_io_result)
  );
  _ x212_1 ( // @[Math.scala 720:24:@4855.4]
    .io_b(x212_1_io_b),
    .io_result(x212_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4868.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@4877.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@4888.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x198_fifoinpacked_0_full; // @[sm_x216_inr_Foreach.scala 62:18:@4774.4]
  assign _T_328 = ~ io_in_x198_fifoinpacked_0_active_0_out; // @[sm_x216_inr_Foreach.scala 62:55:@4775.4]
  assign b203_number = __io_result; // @[Math.scala 723:22:@4754.4 Math.scala 724:14:@4755.4]
  assign _GEN_0 = {{11'd0}, b203_number}; // @[Math.scala 461:32:@4779.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@4779.4]
  assign _GEN_1 = {{7'd0}, b203_number}; // @[Math.scala 461:32:@4784.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@4784.4]
  assign x209_sum_number = x209_sum_1_io_result; // @[Math.scala 154:22:@4825.4 Math.scala 155:14:@4826.4]
  assign _GEN_2 = {{2'd0}, x209_sum_number}; // @[Math.scala 461:32:@4830.4]
  assign _T_353 = _GEN_2 << 2; // @[Math.scala 461:32:@4830.4]
  assign x392_sum_number = x392_sum_1_io_result; // @[Math.scala 154:22:@4840.4 Math.scala 155:14:@4841.4]
  assign _T_364 = $signed(x392_sum_number); // @[Math.scala 406:49:@4847.4]
  assign _T_366 = $signed(_T_364) & $signed(32'shff); // @[Math.scala 406:56:@4849.4]
  assign _T_367 = $signed(_T_366); // @[Math.scala 406:56:@4850.4]
  assign _T_385 = ~ io_sigsIn_break; // @[sm_x216_inr_Foreach.scala 93:131:@4885.4]
  assign _T_389 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4893.4 package.scala 96:25:@4894.4]
  assign _T_391 = io_rr ? _T_389 : 1'h0; // @[implicits.scala 55:10:@4895.4]
  assign _T_392 = _T_385 & _T_391; // @[sm_x216_inr_Foreach.scala 93:148:@4896.4]
  assign _T_394 = _T_392 & _T_385; // @[sm_x216_inr_Foreach.scala 93:236:@4898.4]
  assign _T_395 = _T_394 & io_sigsIn_backpressure; // @[sm_x216_inr_Foreach.scala 93:255:@4899.4]
  assign x478_b205_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4873.4 package.scala 96:25:@4874.4]
  assign _T_398 = _T_395 & x478_b205_D4; // @[sm_x216_inr_Foreach.scala 93:291:@4901.4]
  assign x479_b206_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4882.4 package.scala 96:25:@4883.4]
  assign io_in_x198_fifoinpacked_0_wPort_0_en_0 = _T_398 & x479_b206_D4; // @[MemInterfaceType.scala 93:57:@4905.4]
  assign io_in_x198_fifoinpacked_0_active_0_in = x478_b205_D4 & x479_b206_D4; // @[MemInterfaceType.scala 147:18:@4908.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4752.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@4764.4]
  assign x390_sub_1_clock = clock; // @[:@4789.4]
  assign x390_sub_1_reset = reset; // @[:@4790.4]
  assign x390_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@4791.4]
  assign x390_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@4792.4]
  assign x390_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@4793.4]
  assign RetimeWrapper_clock = clock; // @[:@4799.4]
  assign RetimeWrapper_reset = reset; // @[:@4800.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4802.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@4801.4]
  assign x208_sum_1_clock = clock; // @[:@4808.4]
  assign x208_sum_1_reset = reset; // @[:@4809.4]
  assign x208_sum_1_io_a = x390_sub_1_io_result; // @[Math.scala 151:17:@4810.4]
  assign x208_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@4811.4]
  assign x208_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4812.4]
  assign x209_sum_1_clock = clock; // @[:@4820.4]
  assign x209_sum_1_reset = reset; // @[:@4821.4]
  assign x209_sum_1_io_a = x208_sum_1_io_result; // @[Math.scala 151:17:@4822.4]
  assign x209_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@4823.4]
  assign x209_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4824.4]
  assign x392_sum_1_clock = clock; // @[:@4835.4]
  assign x392_sum_1_reset = reset; // @[:@4836.4]
  assign x392_sum_1_io_a = _T_353[31:0]; // @[Math.scala 151:17:@4837.4]
  assign x392_sum_1_io_b = x209_sum_1_io_result; // @[Math.scala 152:17:@4838.4]
  assign x392_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4839.4]
  assign x212_1_io_b = $unsigned(_T_367); // @[Math.scala 721:17:@4858.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4869.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4870.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4872.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4871.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4878.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4879.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4881.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@4880.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4889.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4890.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4892.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4891.4]
endmodule
module RetimeWrapper_42( // @[:@6026.2]
  input   clock, // @[:@6027.4]
  input   reset, // @[:@6028.4]
  input   io_flow, // @[:@6029.4]
  input   io_in, // @[:@6029.4]
  output  io_out // @[:@6029.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(76)) sr ( // @[RetimeShiftRegister.scala 15:20:@6031.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6044.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6043.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6042.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6041.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6040.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6038.4]
endmodule
module RetimeWrapper_46( // @[:@6154.2]
  input   clock, // @[:@6155.4]
  input   reset, // @[:@6156.4]
  input   io_flow, // @[:@6157.4]
  input   io_in, // @[:@6157.4]
  output  io_out // @[:@6157.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(75)) sr ( // @[RetimeShiftRegister.scala 15:20:@6159.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6172.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6171.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6170.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6169.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6168.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6166.4]
endmodule
module x339_inr_Foreach_SAMPLER_BOX_sm( // @[:@6174.2]
  input   clock, // @[:@6175.4]
  input   reset, // @[:@6176.4]
  input   io_enable, // @[:@6177.4]
  output  io_done, // @[:@6177.4]
  output  io_doneLatch, // @[:@6177.4]
  input   io_ctrDone, // @[:@6177.4]
  output  io_datapathEn, // @[:@6177.4]
  output  io_ctrInc, // @[:@6177.4]
  output  io_ctrRst, // @[:@6177.4]
  input   io_parentAck, // @[:@6177.4]
  input   io_backpressure, // @[:@6177.4]
  input   io_break // @[:@6177.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6179.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6179.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6182.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6182.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6274.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6187.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6188.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6189.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6190.4]
  wire  _T_100; // @[package.scala 100:49:@6207.4]
  reg  _T_103; // @[package.scala 48:56:@6208.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6221.4 package.scala 96:25:@6222.4]
  wire  _T_110; // @[package.scala 100:49:@6223.4]
  reg  _T_113; // @[package.scala 48:56:@6224.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6226.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6231.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6232.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6235.4]
  wire  _T_124; // @[package.scala 96:25:@6243.4 package.scala 96:25:@6244.4]
  wire  _T_126; // @[package.scala 100:49:@6245.4]
  reg  _T_129; // @[package.scala 48:56:@6246.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6268.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6270.4]
  reg  _T_153; // @[package.scala 48:56:@6271.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6279.4 package.scala 96:25:@6280.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6281.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6282.4]
  SRFF active ( // @[Controllers.scala 261:22:@6179.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6182.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_42 RetimeWrapper ( // @[package.scala 93:22:@6216.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_1 ( // @[package.scala 93:22:@6238.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6250.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6258.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_4 ( // @[package.scala 93:22:@6274.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6187.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6188.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6189.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6190.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6207.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6221.4 package.scala 96:25:@6222.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6223.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6226.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6231.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6232.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6235.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6243.4 package.scala 96:25:@6244.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6245.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6270.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6279.4 package.scala 96:25:@6280.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6281.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6282.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6249.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6284.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6234.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6237.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6229.4]
  assign active_clock = clock; // @[:@6180.4]
  assign active_reset = reset; // @[:@6181.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6192.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6196.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6197.4]
  assign done_clock = clock; // @[:@6183.4]
  assign done_reset = reset; // @[:@6184.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6212.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6205.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6206.4]
  assign RetimeWrapper_clock = clock; // @[:@6217.4]
  assign RetimeWrapper_reset = reset; // @[:@6218.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6220.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6219.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6239.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6240.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6242.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6241.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6251.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6252.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6254.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6253.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6259.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6260.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6262.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6261.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6275.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6276.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6278.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6277.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SRAM_1( // @[:@6511.2]
  input         clock, // @[:@6512.4]
  input         reset, // @[:@6513.4]
  input  [9:0]  io_raddr, // @[:@6514.4]
  input         io_wen, // @[:@6514.4]
  input  [9:0]  io_waddr, // @[:@6514.4]
  input  [31:0] io_wdata, // @[:@6514.4]
  output [31:0] io_rdata, // @[:@6514.4]
  input         io_backpressure // @[:@6514.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6516.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6516.4]
  wire [9:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6516.4]
  wire [9:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6516.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6534.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6535.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6536.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6538.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(640), .AWIDTH(10)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6516.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6534.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6535.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6543.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6530.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6531.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6528.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6533.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6532.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6529.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6527.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6526.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_51( // @[:@6557.2]
  input        clock, // @[:@6558.4]
  input        reset, // @[:@6559.4]
  input        io_flow, // @[:@6560.4]
  input  [9:0] io_in, // @[:@6560.4]
  output [9:0] io_out // @[:@6560.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6562.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6575.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6574.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@6573.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6572.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6571.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6569.4]
endmodule
module Mem1D_5( // @[:@6577.2]
  input         clock, // @[:@6578.4]
  input         reset, // @[:@6579.4]
  input  [9:0]  io_r_ofs_0, // @[:@6580.4]
  input         io_r_backpressure, // @[:@6580.4]
  input  [9:0]  io_w_ofs_0, // @[:@6580.4]
  input  [31:0] io_w_data_0, // @[:@6580.4]
  input         io_w_en_0, // @[:@6580.4]
  output [31:0] io_output // @[:@6580.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [9:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [9:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6587.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6587.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6587.4]
  wire [9:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6587.4]
  wire [9:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6587.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@6582.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@6584.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_51 RetimeWrapper ( // @[package.scala 93:22:@6587.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 10'h280; // @[MemPrimitives.scala 702:32:@6582.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@6600.4]
  assign SRAM_clock = clock; // @[:@6585.4]
  assign SRAM_reset = reset; // @[:@6586.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@6594.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@6597.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@6595.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@6598.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@6599.4]
  assign RetimeWrapper_clock = clock; // @[:@6588.4]
  assign RetimeWrapper_reset = reset; // @[:@6589.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@6591.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@6590.4]
endmodule
module StickySelects_1( // @[:@7779.2]
  input   clock, // @[:@7780.4]
  input   reset, // @[:@7781.4]
  input   io_ins_0, // @[:@7782.4]
  input   io_ins_1, // @[:@7782.4]
  input   io_ins_2, // @[:@7782.4]
  input   io_ins_3, // @[:@7782.4]
  input   io_ins_4, // @[:@7782.4]
  input   io_ins_5, // @[:@7782.4]
  input   io_ins_6, // @[:@7782.4]
  input   io_ins_7, // @[:@7782.4]
  input   io_ins_8, // @[:@7782.4]
  output  io_outs_0, // @[:@7782.4]
  output  io_outs_1, // @[:@7782.4]
  output  io_outs_2, // @[:@7782.4]
  output  io_outs_3, // @[:@7782.4]
  output  io_outs_4, // @[:@7782.4]
  output  io_outs_5, // @[:@7782.4]
  output  io_outs_6, // @[:@7782.4]
  output  io_outs_7, // @[:@7782.4]
  output  io_outs_8 // @[:@7782.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@7784.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@7785.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@7786.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@7787.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@7788.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@7789.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@7790.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@7791.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@7792.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@7793.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@7794.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@7795.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@7796.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@7797.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@7798.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@7799.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@7800.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@7801.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@7803.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@7804.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@7805.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@7806.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@7807.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@7808.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@7809.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@7810.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@7811.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@7813.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@7814.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@7815.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@7816.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@7817.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@7818.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@7819.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@7820.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@7821.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@7824.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@7825.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@7826.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@7827.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@7828.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@7829.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@7830.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@7831.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@7835.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@7836.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@7837.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@7838.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@7839.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@7840.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@7841.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@7846.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@7847.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@7848.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@7849.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@7850.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@7851.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@7857.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@7858.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@7859.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@7860.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@7861.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@7868.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@7869.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@7870.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@7871.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@7879.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@7880.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@7881.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@7793.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@7794.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@7795.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@7796.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@7797.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@7798.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@7799.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@7800.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@7801.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@7803.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@7804.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@7805.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@7806.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@7807.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@7808.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@7809.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@7810.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@7811.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@7813.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@7814.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@7815.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@7816.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@7817.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@7818.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@7819.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@7820.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@7821.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@7824.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@7825.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@7826.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@7827.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@7828.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@7829.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@7830.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@7831.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@7835.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@7836.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@7837.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@7838.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@7839.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@7840.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@7841.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@7846.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@7847.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@7848.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@7849.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@7850.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@7851.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@7857.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@7858.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@7859.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@7860.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@7861.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@7868.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@7869.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@7870.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@7871.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@7879.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@7880.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@7881.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@7883.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@7884.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@7885.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@7886.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@7887.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@7888.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@7889.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@7890.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@7891.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x227_lb_0( // @[:@12603.2]
  input         clock, // @[:@12604.4]
  input         reset, // @[:@12605.4]
  input  [1:0]  io_rPort_8_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_8_ofs_0, // @[:@12606.4]
  input         io_rPort_8_en_0, // @[:@12606.4]
  input         io_rPort_8_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_8_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_7_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_7_ofs_0, // @[:@12606.4]
  input         io_rPort_7_en_0, // @[:@12606.4]
  input         io_rPort_7_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_7_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_6_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_6_ofs_0, // @[:@12606.4]
  input         io_rPort_6_en_0, // @[:@12606.4]
  input         io_rPort_6_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_6_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_5_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_5_ofs_0, // @[:@12606.4]
  input         io_rPort_5_en_0, // @[:@12606.4]
  input         io_rPort_5_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_5_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_4_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_4_ofs_0, // @[:@12606.4]
  input         io_rPort_4_en_0, // @[:@12606.4]
  input         io_rPort_4_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_4_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_3_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_3_ofs_0, // @[:@12606.4]
  input         io_rPort_3_en_0, // @[:@12606.4]
  input         io_rPort_3_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_3_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_2_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_2_ofs_0, // @[:@12606.4]
  input         io_rPort_2_en_0, // @[:@12606.4]
  input         io_rPort_2_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_2_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_1_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_1_ofs_0, // @[:@12606.4]
  input         io_rPort_1_en_0, // @[:@12606.4]
  input         io_rPort_1_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_1_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_0_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_0_ofs_0, // @[:@12606.4]
  input         io_rPort_0_en_0, // @[:@12606.4]
  input         io_rPort_0_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_0_output_0, // @[:@12606.4]
  input  [1:0]  io_wPort_0_banks_1, // @[:@12606.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12606.4]
  input  [9:0]  io_wPort_0_ofs_0, // @[:@12606.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12606.4]
  input         io_wPort_0_en_0 // @[:@12606.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [9:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [9:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [9:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [9:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [9:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [9:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [9:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [9:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [9:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [9:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [9:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [9:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [9:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [9:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [9:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [9:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [9:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [9:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [9:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [9:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [9:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [9:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [9:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [9:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@15352.4]
  wire  _T_316; // @[MemPrimitives.scala 82:210:@12863.4]
  wire  _T_318; // @[MemPrimitives.scala 82:210:@12864.4]
  wire  _T_319; // @[MemPrimitives.scala 82:228:@12865.4]
  wire  _T_320; // @[MemPrimitives.scala 83:102:@12866.4]
  wire [42:0] _T_322; // @[Cat.scala 30:58:@12868.4]
  wire  _T_329; // @[MemPrimitives.scala 82:210:@12876.4]
  wire  _T_330; // @[MemPrimitives.scala 82:228:@12877.4]
  wire  _T_331; // @[MemPrimitives.scala 83:102:@12878.4]
  wire [42:0] _T_333; // @[Cat.scala 30:58:@12880.4]
  wire  _T_340; // @[MemPrimitives.scala 82:210:@12888.4]
  wire  _T_341; // @[MemPrimitives.scala 82:228:@12889.4]
  wire  _T_342; // @[MemPrimitives.scala 83:102:@12890.4]
  wire [42:0] _T_344; // @[Cat.scala 30:58:@12892.4]
  wire  _T_349; // @[MemPrimitives.scala 82:210:@12899.4]
  wire  _T_352; // @[MemPrimitives.scala 82:228:@12901.4]
  wire  _T_353; // @[MemPrimitives.scala 83:102:@12902.4]
  wire [42:0] _T_355; // @[Cat.scala 30:58:@12904.4]
  wire  _T_363; // @[MemPrimitives.scala 82:228:@12913.4]
  wire  _T_364; // @[MemPrimitives.scala 83:102:@12914.4]
  wire [42:0] _T_366; // @[Cat.scala 30:58:@12916.4]
  wire  _T_374; // @[MemPrimitives.scala 82:228:@12925.4]
  wire  _T_375; // @[MemPrimitives.scala 83:102:@12926.4]
  wire [42:0] _T_377; // @[Cat.scala 30:58:@12928.4]
  wire  _T_382; // @[MemPrimitives.scala 82:210:@12935.4]
  wire  _T_385; // @[MemPrimitives.scala 82:228:@12937.4]
  wire  _T_386; // @[MemPrimitives.scala 83:102:@12938.4]
  wire [42:0] _T_388; // @[Cat.scala 30:58:@12940.4]
  wire  _T_396; // @[MemPrimitives.scala 82:228:@12949.4]
  wire  _T_397; // @[MemPrimitives.scala 83:102:@12950.4]
  wire [42:0] _T_399; // @[Cat.scala 30:58:@12952.4]
  wire  _T_407; // @[MemPrimitives.scala 82:228:@12961.4]
  wire  _T_408; // @[MemPrimitives.scala 83:102:@12962.4]
  wire [42:0] _T_410; // @[Cat.scala 30:58:@12964.4]
  wire  _T_415; // @[MemPrimitives.scala 82:210:@12971.4]
  wire  _T_418; // @[MemPrimitives.scala 82:228:@12973.4]
  wire  _T_419; // @[MemPrimitives.scala 83:102:@12974.4]
  wire [42:0] _T_421; // @[Cat.scala 30:58:@12976.4]
  wire  _T_429; // @[MemPrimitives.scala 82:228:@12985.4]
  wire  _T_430; // @[MemPrimitives.scala 83:102:@12986.4]
  wire [42:0] _T_432; // @[Cat.scala 30:58:@12988.4]
  wire  _T_440; // @[MemPrimitives.scala 82:228:@12997.4]
  wire  _T_441; // @[MemPrimitives.scala 83:102:@12998.4]
  wire [42:0] _T_443; // @[Cat.scala 30:58:@13000.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@13007.4]
  wire  _T_450; // @[MemPrimitives.scala 110:210:@13008.4]
  wire  _T_451; // @[MemPrimitives.scala 110:228:@13009.4]
  wire  _T_454; // @[MemPrimitives.scala 110:210:@13011.4]
  wire  _T_456; // @[MemPrimitives.scala 110:210:@13012.4]
  wire  _T_457; // @[MemPrimitives.scala 110:228:@13013.4]
  wire  _T_460; // @[MemPrimitives.scala 110:210:@13015.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@13016.4]
  wire  _T_463; // @[MemPrimitives.scala 110:228:@13017.4]
  wire  _T_466; // @[MemPrimitives.scala 110:210:@13019.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@13020.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@13021.4]
  wire  _T_472; // @[MemPrimitives.scala 110:210:@13023.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@13024.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@13025.4]
  wire  _T_478; // @[MemPrimitives.scala 110:210:@13027.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@13028.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@13029.4]
  wire  _T_484; // @[MemPrimitives.scala 110:210:@13031.4]
  wire  _T_486; // @[MemPrimitives.scala 110:210:@13032.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@13033.4]
  wire  _T_490; // @[MemPrimitives.scala 110:210:@13035.4]
  wire  _T_492; // @[MemPrimitives.scala 110:210:@13036.4]
  wire  _T_493; // @[MemPrimitives.scala 110:228:@13037.4]
  wire  _T_496; // @[MemPrimitives.scala 110:210:@13039.4]
  wire  _T_498; // @[MemPrimitives.scala 110:210:@13040.4]
  wire  _T_499; // @[MemPrimitives.scala 110:228:@13041.4]
  wire  _T_501; // @[MemPrimitives.scala 126:35:@13055.4]
  wire  _T_502; // @[MemPrimitives.scala 126:35:@13056.4]
  wire  _T_503; // @[MemPrimitives.scala 126:35:@13057.4]
  wire  _T_504; // @[MemPrimitives.scala 126:35:@13058.4]
  wire  _T_505; // @[MemPrimitives.scala 126:35:@13059.4]
  wire  _T_506; // @[MemPrimitives.scala 126:35:@13060.4]
  wire  _T_507; // @[MemPrimitives.scala 126:35:@13061.4]
  wire  _T_508; // @[MemPrimitives.scala 126:35:@13062.4]
  wire  _T_509; // @[MemPrimitives.scala 126:35:@13063.4]
  wire [11:0] _T_511; // @[Cat.scala 30:58:@13065.4]
  wire [11:0] _T_513; // @[Cat.scala 30:58:@13067.4]
  wire [11:0] _T_515; // @[Cat.scala 30:58:@13069.4]
  wire [11:0] _T_517; // @[Cat.scala 30:58:@13071.4]
  wire [11:0] _T_519; // @[Cat.scala 30:58:@13073.4]
  wire [11:0] _T_521; // @[Cat.scala 30:58:@13075.4]
  wire [11:0] _T_523; // @[Cat.scala 30:58:@13077.4]
  wire [11:0] _T_525; // @[Cat.scala 30:58:@13079.4]
  wire [11:0] _T_527; // @[Cat.scala 30:58:@13081.4]
  wire [11:0] _T_528; // @[Mux.scala 31:69:@13082.4]
  wire [11:0] _T_529; // @[Mux.scala 31:69:@13083.4]
  wire [11:0] _T_530; // @[Mux.scala 31:69:@13084.4]
  wire [11:0] _T_531; // @[Mux.scala 31:69:@13085.4]
  wire [11:0] _T_532; // @[Mux.scala 31:69:@13086.4]
  wire [11:0] _T_533; // @[Mux.scala 31:69:@13087.4]
  wire [11:0] _T_534; // @[Mux.scala 31:69:@13088.4]
  wire [11:0] _T_535; // @[Mux.scala 31:69:@13089.4]
  wire  _T_542; // @[MemPrimitives.scala 110:210:@13097.4]
  wire  _T_543; // @[MemPrimitives.scala 110:228:@13098.4]
  wire  _T_548; // @[MemPrimitives.scala 110:210:@13101.4]
  wire  _T_549; // @[MemPrimitives.scala 110:228:@13102.4]
  wire  _T_554; // @[MemPrimitives.scala 110:210:@13105.4]
  wire  _T_555; // @[MemPrimitives.scala 110:228:@13106.4]
  wire  _T_560; // @[MemPrimitives.scala 110:210:@13109.4]
  wire  _T_561; // @[MemPrimitives.scala 110:228:@13110.4]
  wire  _T_566; // @[MemPrimitives.scala 110:210:@13113.4]
  wire  _T_567; // @[MemPrimitives.scala 110:228:@13114.4]
  wire  _T_572; // @[MemPrimitives.scala 110:210:@13117.4]
  wire  _T_573; // @[MemPrimitives.scala 110:228:@13118.4]
  wire  _T_578; // @[MemPrimitives.scala 110:210:@13121.4]
  wire  _T_579; // @[MemPrimitives.scala 110:228:@13122.4]
  wire  _T_584; // @[MemPrimitives.scala 110:210:@13125.4]
  wire  _T_585; // @[MemPrimitives.scala 110:228:@13126.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@13129.4]
  wire  _T_591; // @[MemPrimitives.scala 110:228:@13130.4]
  wire  _T_593; // @[MemPrimitives.scala 126:35:@13144.4]
  wire  _T_594; // @[MemPrimitives.scala 126:35:@13145.4]
  wire  _T_595; // @[MemPrimitives.scala 126:35:@13146.4]
  wire  _T_596; // @[MemPrimitives.scala 126:35:@13147.4]
  wire  _T_597; // @[MemPrimitives.scala 126:35:@13148.4]
  wire  _T_598; // @[MemPrimitives.scala 126:35:@13149.4]
  wire  _T_599; // @[MemPrimitives.scala 126:35:@13150.4]
  wire  _T_600; // @[MemPrimitives.scala 126:35:@13151.4]
  wire  _T_601; // @[MemPrimitives.scala 126:35:@13152.4]
  wire [11:0] _T_603; // @[Cat.scala 30:58:@13154.4]
  wire [11:0] _T_605; // @[Cat.scala 30:58:@13156.4]
  wire [11:0] _T_607; // @[Cat.scala 30:58:@13158.4]
  wire [11:0] _T_609; // @[Cat.scala 30:58:@13160.4]
  wire [11:0] _T_611; // @[Cat.scala 30:58:@13162.4]
  wire [11:0] _T_613; // @[Cat.scala 30:58:@13164.4]
  wire [11:0] _T_615; // @[Cat.scala 30:58:@13166.4]
  wire [11:0] _T_617; // @[Cat.scala 30:58:@13168.4]
  wire [11:0] _T_619; // @[Cat.scala 30:58:@13170.4]
  wire [11:0] _T_620; // @[Mux.scala 31:69:@13171.4]
  wire [11:0] _T_621; // @[Mux.scala 31:69:@13172.4]
  wire [11:0] _T_622; // @[Mux.scala 31:69:@13173.4]
  wire [11:0] _T_623; // @[Mux.scala 31:69:@13174.4]
  wire [11:0] _T_624; // @[Mux.scala 31:69:@13175.4]
  wire [11:0] _T_625; // @[Mux.scala 31:69:@13176.4]
  wire [11:0] _T_626; // @[Mux.scala 31:69:@13177.4]
  wire [11:0] _T_627; // @[Mux.scala 31:69:@13178.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@13186.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@13187.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13190.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@13191.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13194.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13195.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13198.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13199.4]
  wire  _T_658; // @[MemPrimitives.scala 110:210:@13202.4]
  wire  _T_659; // @[MemPrimitives.scala 110:228:@13203.4]
  wire  _T_664; // @[MemPrimitives.scala 110:210:@13206.4]
  wire  _T_665; // @[MemPrimitives.scala 110:228:@13207.4]
  wire  _T_670; // @[MemPrimitives.scala 110:210:@13210.4]
  wire  _T_671; // @[MemPrimitives.scala 110:228:@13211.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@13214.4]
  wire  _T_677; // @[MemPrimitives.scala 110:228:@13215.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13218.4]
  wire  _T_683; // @[MemPrimitives.scala 110:228:@13219.4]
  wire  _T_685; // @[MemPrimitives.scala 126:35:@13233.4]
  wire  _T_686; // @[MemPrimitives.scala 126:35:@13234.4]
  wire  _T_687; // @[MemPrimitives.scala 126:35:@13235.4]
  wire  _T_688; // @[MemPrimitives.scala 126:35:@13236.4]
  wire  _T_689; // @[MemPrimitives.scala 126:35:@13237.4]
  wire  _T_690; // @[MemPrimitives.scala 126:35:@13238.4]
  wire  _T_691; // @[MemPrimitives.scala 126:35:@13239.4]
  wire  _T_692; // @[MemPrimitives.scala 126:35:@13240.4]
  wire  _T_693; // @[MemPrimitives.scala 126:35:@13241.4]
  wire [11:0] _T_695; // @[Cat.scala 30:58:@13243.4]
  wire [11:0] _T_697; // @[Cat.scala 30:58:@13245.4]
  wire [11:0] _T_699; // @[Cat.scala 30:58:@13247.4]
  wire [11:0] _T_701; // @[Cat.scala 30:58:@13249.4]
  wire [11:0] _T_703; // @[Cat.scala 30:58:@13251.4]
  wire [11:0] _T_705; // @[Cat.scala 30:58:@13253.4]
  wire [11:0] _T_707; // @[Cat.scala 30:58:@13255.4]
  wire [11:0] _T_709; // @[Cat.scala 30:58:@13257.4]
  wire [11:0] _T_711; // @[Cat.scala 30:58:@13259.4]
  wire [11:0] _T_712; // @[Mux.scala 31:69:@13260.4]
  wire [11:0] _T_713; // @[Mux.scala 31:69:@13261.4]
  wire [11:0] _T_714; // @[Mux.scala 31:69:@13262.4]
  wire [11:0] _T_715; // @[Mux.scala 31:69:@13263.4]
  wire [11:0] _T_716; // @[Mux.scala 31:69:@13264.4]
  wire [11:0] _T_717; // @[Mux.scala 31:69:@13265.4]
  wire [11:0] _T_718; // @[Mux.scala 31:69:@13266.4]
  wire [11:0] _T_719; // @[Mux.scala 31:69:@13267.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@13274.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@13276.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@13278.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@13280.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@13282.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@13284.4]
  wire  _T_742; // @[MemPrimitives.scala 110:210:@13286.4]
  wire  _T_745; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_748; // @[MemPrimitives.scala 110:210:@13290.4]
  wire  _T_751; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_754; // @[MemPrimitives.scala 110:210:@13294.4]
  wire  _T_757; // @[MemPrimitives.scala 110:228:@13296.4]
  wire  _T_760; // @[MemPrimitives.scala 110:210:@13298.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@13300.4]
  wire  _T_766; // @[MemPrimitives.scala 110:210:@13302.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@13304.4]
  wire  _T_772; // @[MemPrimitives.scala 110:210:@13306.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@13308.4]
  wire  _T_777; // @[MemPrimitives.scala 126:35:@13322.4]
  wire  _T_778; // @[MemPrimitives.scala 126:35:@13323.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@13324.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@13325.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@13326.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@13327.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@13328.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@13329.4]
  wire  _T_785; // @[MemPrimitives.scala 126:35:@13330.4]
  wire [11:0] _T_787; // @[Cat.scala 30:58:@13332.4]
  wire [11:0] _T_789; // @[Cat.scala 30:58:@13334.4]
  wire [11:0] _T_791; // @[Cat.scala 30:58:@13336.4]
  wire [11:0] _T_793; // @[Cat.scala 30:58:@13338.4]
  wire [11:0] _T_795; // @[Cat.scala 30:58:@13340.4]
  wire [11:0] _T_797; // @[Cat.scala 30:58:@13342.4]
  wire [11:0] _T_799; // @[Cat.scala 30:58:@13344.4]
  wire [11:0] _T_801; // @[Cat.scala 30:58:@13346.4]
  wire [11:0] _T_803; // @[Cat.scala 30:58:@13348.4]
  wire [11:0] _T_804; // @[Mux.scala 31:69:@13349.4]
  wire [11:0] _T_805; // @[Mux.scala 31:69:@13350.4]
  wire [11:0] _T_806; // @[Mux.scala 31:69:@13351.4]
  wire [11:0] _T_807; // @[Mux.scala 31:69:@13352.4]
  wire [11:0] _T_808; // @[Mux.scala 31:69:@13353.4]
  wire [11:0] _T_809; // @[Mux.scala 31:69:@13354.4]
  wire [11:0] _T_810; // @[Mux.scala 31:69:@13355.4]
  wire [11:0] _T_811; // @[Mux.scala 31:69:@13356.4]
  wire  _T_819; // @[MemPrimitives.scala 110:228:@13365.4]
  wire  _T_825; // @[MemPrimitives.scala 110:228:@13369.4]
  wire  _T_831; // @[MemPrimitives.scala 110:228:@13373.4]
  wire  _T_837; // @[MemPrimitives.scala 110:228:@13377.4]
  wire  _T_843; // @[MemPrimitives.scala 110:228:@13381.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@13385.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@13389.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@13393.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@13397.4]
  wire  _T_869; // @[MemPrimitives.scala 126:35:@13411.4]
  wire  _T_870; // @[MemPrimitives.scala 126:35:@13412.4]
  wire  _T_871; // @[MemPrimitives.scala 126:35:@13413.4]
  wire  _T_872; // @[MemPrimitives.scala 126:35:@13414.4]
  wire  _T_873; // @[MemPrimitives.scala 126:35:@13415.4]
  wire  _T_874; // @[MemPrimitives.scala 126:35:@13416.4]
  wire  _T_875; // @[MemPrimitives.scala 126:35:@13417.4]
  wire  _T_876; // @[MemPrimitives.scala 126:35:@13418.4]
  wire  _T_877; // @[MemPrimitives.scala 126:35:@13419.4]
  wire [11:0] _T_879; // @[Cat.scala 30:58:@13421.4]
  wire [11:0] _T_881; // @[Cat.scala 30:58:@13423.4]
  wire [11:0] _T_883; // @[Cat.scala 30:58:@13425.4]
  wire [11:0] _T_885; // @[Cat.scala 30:58:@13427.4]
  wire [11:0] _T_887; // @[Cat.scala 30:58:@13429.4]
  wire [11:0] _T_889; // @[Cat.scala 30:58:@13431.4]
  wire [11:0] _T_891; // @[Cat.scala 30:58:@13433.4]
  wire [11:0] _T_893; // @[Cat.scala 30:58:@13435.4]
  wire [11:0] _T_895; // @[Cat.scala 30:58:@13437.4]
  wire [11:0] _T_896; // @[Mux.scala 31:69:@13438.4]
  wire [11:0] _T_897; // @[Mux.scala 31:69:@13439.4]
  wire [11:0] _T_898; // @[Mux.scala 31:69:@13440.4]
  wire [11:0] _T_899; // @[Mux.scala 31:69:@13441.4]
  wire [11:0] _T_900; // @[Mux.scala 31:69:@13442.4]
  wire [11:0] _T_901; // @[Mux.scala 31:69:@13443.4]
  wire [11:0] _T_902; // @[Mux.scala 31:69:@13444.4]
  wire [11:0] _T_903; // @[Mux.scala 31:69:@13445.4]
  wire  _T_911; // @[MemPrimitives.scala 110:228:@13454.4]
  wire  _T_917; // @[MemPrimitives.scala 110:228:@13458.4]
  wire  _T_923; // @[MemPrimitives.scala 110:228:@13462.4]
  wire  _T_929; // @[MemPrimitives.scala 110:228:@13466.4]
  wire  _T_935; // @[MemPrimitives.scala 110:228:@13470.4]
  wire  _T_941; // @[MemPrimitives.scala 110:228:@13474.4]
  wire  _T_947; // @[MemPrimitives.scala 110:228:@13478.4]
  wire  _T_953; // @[MemPrimitives.scala 110:228:@13482.4]
  wire  _T_959; // @[MemPrimitives.scala 110:228:@13486.4]
  wire  _T_961; // @[MemPrimitives.scala 126:35:@13500.4]
  wire  _T_962; // @[MemPrimitives.scala 126:35:@13501.4]
  wire  _T_963; // @[MemPrimitives.scala 126:35:@13502.4]
  wire  _T_964; // @[MemPrimitives.scala 126:35:@13503.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13504.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13505.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13506.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13507.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13508.4]
  wire [11:0] _T_971; // @[Cat.scala 30:58:@13510.4]
  wire [11:0] _T_973; // @[Cat.scala 30:58:@13512.4]
  wire [11:0] _T_975; // @[Cat.scala 30:58:@13514.4]
  wire [11:0] _T_977; // @[Cat.scala 30:58:@13516.4]
  wire [11:0] _T_979; // @[Cat.scala 30:58:@13518.4]
  wire [11:0] _T_981; // @[Cat.scala 30:58:@13520.4]
  wire [11:0] _T_983; // @[Cat.scala 30:58:@13522.4]
  wire [11:0] _T_985; // @[Cat.scala 30:58:@13524.4]
  wire [11:0] _T_987; // @[Cat.scala 30:58:@13526.4]
  wire [11:0] _T_988; // @[Mux.scala 31:69:@13527.4]
  wire [11:0] _T_989; // @[Mux.scala 31:69:@13528.4]
  wire [11:0] _T_990; // @[Mux.scala 31:69:@13529.4]
  wire [11:0] _T_991; // @[Mux.scala 31:69:@13530.4]
  wire [11:0] _T_992; // @[Mux.scala 31:69:@13531.4]
  wire [11:0] _T_993; // @[Mux.scala 31:69:@13532.4]
  wire [11:0] _T_994; // @[Mux.scala 31:69:@13533.4]
  wire [11:0] _T_995; // @[Mux.scala 31:69:@13534.4]
  wire  _T_1000; // @[MemPrimitives.scala 110:210:@13541.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@13543.4]
  wire  _T_1006; // @[MemPrimitives.scala 110:210:@13545.4]
  wire  _T_1009; // @[MemPrimitives.scala 110:228:@13547.4]
  wire  _T_1012; // @[MemPrimitives.scala 110:210:@13549.4]
  wire  _T_1015; // @[MemPrimitives.scala 110:228:@13551.4]
  wire  _T_1018; // @[MemPrimitives.scala 110:210:@13553.4]
  wire  _T_1021; // @[MemPrimitives.scala 110:228:@13555.4]
  wire  _T_1024; // @[MemPrimitives.scala 110:210:@13557.4]
  wire  _T_1027; // @[MemPrimitives.scala 110:228:@13559.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@13561.4]
  wire  _T_1033; // @[MemPrimitives.scala 110:228:@13563.4]
  wire  _T_1036; // @[MemPrimitives.scala 110:210:@13565.4]
  wire  _T_1039; // @[MemPrimitives.scala 110:228:@13567.4]
  wire  _T_1042; // @[MemPrimitives.scala 110:210:@13569.4]
  wire  _T_1045; // @[MemPrimitives.scala 110:228:@13571.4]
  wire  _T_1048; // @[MemPrimitives.scala 110:210:@13573.4]
  wire  _T_1051; // @[MemPrimitives.scala 110:228:@13575.4]
  wire  _T_1053; // @[MemPrimitives.scala 126:35:@13589.4]
  wire  _T_1054; // @[MemPrimitives.scala 126:35:@13590.4]
  wire  _T_1055; // @[MemPrimitives.scala 126:35:@13591.4]
  wire  _T_1056; // @[MemPrimitives.scala 126:35:@13592.4]
  wire  _T_1057; // @[MemPrimitives.scala 126:35:@13593.4]
  wire  _T_1058; // @[MemPrimitives.scala 126:35:@13594.4]
  wire  _T_1059; // @[MemPrimitives.scala 126:35:@13595.4]
  wire  _T_1060; // @[MemPrimitives.scala 126:35:@13596.4]
  wire  _T_1061; // @[MemPrimitives.scala 126:35:@13597.4]
  wire [11:0] _T_1063; // @[Cat.scala 30:58:@13599.4]
  wire [11:0] _T_1065; // @[Cat.scala 30:58:@13601.4]
  wire [11:0] _T_1067; // @[Cat.scala 30:58:@13603.4]
  wire [11:0] _T_1069; // @[Cat.scala 30:58:@13605.4]
  wire [11:0] _T_1071; // @[Cat.scala 30:58:@13607.4]
  wire [11:0] _T_1073; // @[Cat.scala 30:58:@13609.4]
  wire [11:0] _T_1075; // @[Cat.scala 30:58:@13611.4]
  wire [11:0] _T_1077; // @[Cat.scala 30:58:@13613.4]
  wire [11:0] _T_1079; // @[Cat.scala 30:58:@13615.4]
  wire [11:0] _T_1080; // @[Mux.scala 31:69:@13616.4]
  wire [11:0] _T_1081; // @[Mux.scala 31:69:@13617.4]
  wire [11:0] _T_1082; // @[Mux.scala 31:69:@13618.4]
  wire [11:0] _T_1083; // @[Mux.scala 31:69:@13619.4]
  wire [11:0] _T_1084; // @[Mux.scala 31:69:@13620.4]
  wire [11:0] _T_1085; // @[Mux.scala 31:69:@13621.4]
  wire [11:0] _T_1086; // @[Mux.scala 31:69:@13622.4]
  wire [11:0] _T_1087; // @[Mux.scala 31:69:@13623.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@13632.4]
  wire  _T_1101; // @[MemPrimitives.scala 110:228:@13636.4]
  wire  _T_1107; // @[MemPrimitives.scala 110:228:@13640.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:228:@13644.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13648.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13652.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13656.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13660.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13664.4]
  wire  _T_1145; // @[MemPrimitives.scala 126:35:@13678.4]
  wire  _T_1146; // @[MemPrimitives.scala 126:35:@13679.4]
  wire  _T_1147; // @[MemPrimitives.scala 126:35:@13680.4]
  wire  _T_1148; // @[MemPrimitives.scala 126:35:@13681.4]
  wire  _T_1149; // @[MemPrimitives.scala 126:35:@13682.4]
  wire  _T_1150; // @[MemPrimitives.scala 126:35:@13683.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13684.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13685.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13686.4]
  wire [11:0] _T_1155; // @[Cat.scala 30:58:@13688.4]
  wire [11:0] _T_1157; // @[Cat.scala 30:58:@13690.4]
  wire [11:0] _T_1159; // @[Cat.scala 30:58:@13692.4]
  wire [11:0] _T_1161; // @[Cat.scala 30:58:@13694.4]
  wire [11:0] _T_1163; // @[Cat.scala 30:58:@13696.4]
  wire [11:0] _T_1165; // @[Cat.scala 30:58:@13698.4]
  wire [11:0] _T_1167; // @[Cat.scala 30:58:@13700.4]
  wire [11:0] _T_1169; // @[Cat.scala 30:58:@13702.4]
  wire [11:0] _T_1171; // @[Cat.scala 30:58:@13704.4]
  wire [11:0] _T_1172; // @[Mux.scala 31:69:@13705.4]
  wire [11:0] _T_1173; // @[Mux.scala 31:69:@13706.4]
  wire [11:0] _T_1174; // @[Mux.scala 31:69:@13707.4]
  wire [11:0] _T_1175; // @[Mux.scala 31:69:@13708.4]
  wire [11:0] _T_1176; // @[Mux.scala 31:69:@13709.4]
  wire [11:0] _T_1177; // @[Mux.scala 31:69:@13710.4]
  wire [11:0] _T_1178; // @[Mux.scala 31:69:@13711.4]
  wire [11:0] _T_1179; // @[Mux.scala 31:69:@13712.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13721.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13725.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13729.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13733.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13737.4]
  wire  _T_1217; // @[MemPrimitives.scala 110:228:@13741.4]
  wire  _T_1223; // @[MemPrimitives.scala 110:228:@13745.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:228:@13749.4]
  wire  _T_1235; // @[MemPrimitives.scala 110:228:@13753.4]
  wire  _T_1237; // @[MemPrimitives.scala 126:35:@13767.4]
  wire  _T_1238; // @[MemPrimitives.scala 126:35:@13768.4]
  wire  _T_1239; // @[MemPrimitives.scala 126:35:@13769.4]
  wire  _T_1240; // @[MemPrimitives.scala 126:35:@13770.4]
  wire  _T_1241; // @[MemPrimitives.scala 126:35:@13771.4]
  wire  _T_1242; // @[MemPrimitives.scala 126:35:@13772.4]
  wire  _T_1243; // @[MemPrimitives.scala 126:35:@13773.4]
  wire  _T_1244; // @[MemPrimitives.scala 126:35:@13774.4]
  wire  _T_1245; // @[MemPrimitives.scala 126:35:@13775.4]
  wire [11:0] _T_1247; // @[Cat.scala 30:58:@13777.4]
  wire [11:0] _T_1249; // @[Cat.scala 30:58:@13779.4]
  wire [11:0] _T_1251; // @[Cat.scala 30:58:@13781.4]
  wire [11:0] _T_1253; // @[Cat.scala 30:58:@13783.4]
  wire [11:0] _T_1255; // @[Cat.scala 30:58:@13785.4]
  wire [11:0] _T_1257; // @[Cat.scala 30:58:@13787.4]
  wire [11:0] _T_1259; // @[Cat.scala 30:58:@13789.4]
  wire [11:0] _T_1261; // @[Cat.scala 30:58:@13791.4]
  wire [11:0] _T_1263; // @[Cat.scala 30:58:@13793.4]
  wire [11:0] _T_1264; // @[Mux.scala 31:69:@13794.4]
  wire [11:0] _T_1265; // @[Mux.scala 31:69:@13795.4]
  wire [11:0] _T_1266; // @[Mux.scala 31:69:@13796.4]
  wire [11:0] _T_1267; // @[Mux.scala 31:69:@13797.4]
  wire [11:0] _T_1268; // @[Mux.scala 31:69:@13798.4]
  wire [11:0] _T_1269; // @[Mux.scala 31:69:@13799.4]
  wire [11:0] _T_1270; // @[Mux.scala 31:69:@13800.4]
  wire [11:0] _T_1271; // @[Mux.scala 31:69:@13801.4]
  wire  _T_1276; // @[MemPrimitives.scala 110:210:@13808.4]
  wire  _T_1279; // @[MemPrimitives.scala 110:228:@13810.4]
  wire  _T_1282; // @[MemPrimitives.scala 110:210:@13812.4]
  wire  _T_1285; // @[MemPrimitives.scala 110:228:@13814.4]
  wire  _T_1288; // @[MemPrimitives.scala 110:210:@13816.4]
  wire  _T_1291; // @[MemPrimitives.scala 110:228:@13818.4]
  wire  _T_1294; // @[MemPrimitives.scala 110:210:@13820.4]
  wire  _T_1297; // @[MemPrimitives.scala 110:228:@13822.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@13824.4]
  wire  _T_1303; // @[MemPrimitives.scala 110:228:@13826.4]
  wire  _T_1306; // @[MemPrimitives.scala 110:210:@13828.4]
  wire  _T_1309; // @[MemPrimitives.scala 110:228:@13830.4]
  wire  _T_1312; // @[MemPrimitives.scala 110:210:@13832.4]
  wire  _T_1315; // @[MemPrimitives.scala 110:228:@13834.4]
  wire  _T_1318; // @[MemPrimitives.scala 110:210:@13836.4]
  wire  _T_1321; // @[MemPrimitives.scala 110:228:@13838.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@13840.4]
  wire  _T_1327; // @[MemPrimitives.scala 110:228:@13842.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@13856.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@13857.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@13858.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@13859.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@13860.4]
  wire  _T_1334; // @[MemPrimitives.scala 126:35:@13861.4]
  wire  _T_1335; // @[MemPrimitives.scala 126:35:@13862.4]
  wire  _T_1336; // @[MemPrimitives.scala 126:35:@13863.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13864.4]
  wire [11:0] _T_1339; // @[Cat.scala 30:58:@13866.4]
  wire [11:0] _T_1341; // @[Cat.scala 30:58:@13868.4]
  wire [11:0] _T_1343; // @[Cat.scala 30:58:@13870.4]
  wire [11:0] _T_1345; // @[Cat.scala 30:58:@13872.4]
  wire [11:0] _T_1347; // @[Cat.scala 30:58:@13874.4]
  wire [11:0] _T_1349; // @[Cat.scala 30:58:@13876.4]
  wire [11:0] _T_1351; // @[Cat.scala 30:58:@13878.4]
  wire [11:0] _T_1353; // @[Cat.scala 30:58:@13880.4]
  wire [11:0] _T_1355; // @[Cat.scala 30:58:@13882.4]
  wire [11:0] _T_1356; // @[Mux.scala 31:69:@13883.4]
  wire [11:0] _T_1357; // @[Mux.scala 31:69:@13884.4]
  wire [11:0] _T_1358; // @[Mux.scala 31:69:@13885.4]
  wire [11:0] _T_1359; // @[Mux.scala 31:69:@13886.4]
  wire [11:0] _T_1360; // @[Mux.scala 31:69:@13887.4]
  wire [11:0] _T_1361; // @[Mux.scala 31:69:@13888.4]
  wire [11:0] _T_1362; // @[Mux.scala 31:69:@13889.4]
  wire [11:0] _T_1363; // @[Mux.scala 31:69:@13890.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@13899.4]
  wire  _T_1377; // @[MemPrimitives.scala 110:228:@13903.4]
  wire  _T_1383; // @[MemPrimitives.scala 110:228:@13907.4]
  wire  _T_1389; // @[MemPrimitives.scala 110:228:@13911.4]
  wire  _T_1395; // @[MemPrimitives.scala 110:228:@13915.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:228:@13919.4]
  wire  _T_1407; // @[MemPrimitives.scala 110:228:@13923.4]
  wire  _T_1413; // @[MemPrimitives.scala 110:228:@13927.4]
  wire  _T_1419; // @[MemPrimitives.scala 110:228:@13931.4]
  wire  _T_1421; // @[MemPrimitives.scala 126:35:@13945.4]
  wire  _T_1422; // @[MemPrimitives.scala 126:35:@13946.4]
  wire  _T_1423; // @[MemPrimitives.scala 126:35:@13947.4]
  wire  _T_1424; // @[MemPrimitives.scala 126:35:@13948.4]
  wire  _T_1425; // @[MemPrimitives.scala 126:35:@13949.4]
  wire  _T_1426; // @[MemPrimitives.scala 126:35:@13950.4]
  wire  _T_1427; // @[MemPrimitives.scala 126:35:@13951.4]
  wire  _T_1428; // @[MemPrimitives.scala 126:35:@13952.4]
  wire  _T_1429; // @[MemPrimitives.scala 126:35:@13953.4]
  wire [11:0] _T_1431; // @[Cat.scala 30:58:@13955.4]
  wire [11:0] _T_1433; // @[Cat.scala 30:58:@13957.4]
  wire [11:0] _T_1435; // @[Cat.scala 30:58:@13959.4]
  wire [11:0] _T_1437; // @[Cat.scala 30:58:@13961.4]
  wire [11:0] _T_1439; // @[Cat.scala 30:58:@13963.4]
  wire [11:0] _T_1441; // @[Cat.scala 30:58:@13965.4]
  wire [11:0] _T_1443; // @[Cat.scala 30:58:@13967.4]
  wire [11:0] _T_1445; // @[Cat.scala 30:58:@13969.4]
  wire [11:0] _T_1447; // @[Cat.scala 30:58:@13971.4]
  wire [11:0] _T_1448; // @[Mux.scala 31:69:@13972.4]
  wire [11:0] _T_1449; // @[Mux.scala 31:69:@13973.4]
  wire [11:0] _T_1450; // @[Mux.scala 31:69:@13974.4]
  wire [11:0] _T_1451; // @[Mux.scala 31:69:@13975.4]
  wire [11:0] _T_1452; // @[Mux.scala 31:69:@13976.4]
  wire [11:0] _T_1453; // @[Mux.scala 31:69:@13977.4]
  wire [11:0] _T_1454; // @[Mux.scala 31:69:@13978.4]
  wire [11:0] _T_1455; // @[Mux.scala 31:69:@13979.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@13988.4]
  wire  _T_1469; // @[MemPrimitives.scala 110:228:@13992.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:228:@13996.4]
  wire  _T_1481; // @[MemPrimitives.scala 110:228:@14000.4]
  wire  _T_1487; // @[MemPrimitives.scala 110:228:@14004.4]
  wire  _T_1493; // @[MemPrimitives.scala 110:228:@14008.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:228:@14012.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:228:@14016.4]
  wire  _T_1511; // @[MemPrimitives.scala 110:228:@14020.4]
  wire  _T_1513; // @[MemPrimitives.scala 126:35:@14034.4]
  wire  _T_1514; // @[MemPrimitives.scala 126:35:@14035.4]
  wire  _T_1515; // @[MemPrimitives.scala 126:35:@14036.4]
  wire  _T_1516; // @[MemPrimitives.scala 126:35:@14037.4]
  wire  _T_1517; // @[MemPrimitives.scala 126:35:@14038.4]
  wire  _T_1518; // @[MemPrimitives.scala 126:35:@14039.4]
  wire  _T_1519; // @[MemPrimitives.scala 126:35:@14040.4]
  wire  _T_1520; // @[MemPrimitives.scala 126:35:@14041.4]
  wire  _T_1521; // @[MemPrimitives.scala 126:35:@14042.4]
  wire [11:0] _T_1523; // @[Cat.scala 30:58:@14044.4]
  wire [11:0] _T_1525; // @[Cat.scala 30:58:@14046.4]
  wire [11:0] _T_1527; // @[Cat.scala 30:58:@14048.4]
  wire [11:0] _T_1529; // @[Cat.scala 30:58:@14050.4]
  wire [11:0] _T_1531; // @[Cat.scala 30:58:@14052.4]
  wire [11:0] _T_1533; // @[Cat.scala 30:58:@14054.4]
  wire [11:0] _T_1535; // @[Cat.scala 30:58:@14056.4]
  wire [11:0] _T_1537; // @[Cat.scala 30:58:@14058.4]
  wire [11:0] _T_1539; // @[Cat.scala 30:58:@14060.4]
  wire [11:0] _T_1540; // @[Mux.scala 31:69:@14061.4]
  wire [11:0] _T_1541; // @[Mux.scala 31:69:@14062.4]
  wire [11:0] _T_1542; // @[Mux.scala 31:69:@14063.4]
  wire [11:0] _T_1543; // @[Mux.scala 31:69:@14064.4]
  wire [11:0] _T_1544; // @[Mux.scala 31:69:@14065.4]
  wire [11:0] _T_1545; // @[Mux.scala 31:69:@14066.4]
  wire [11:0] _T_1546; // @[Mux.scala 31:69:@14067.4]
  wire [11:0] _T_1547; // @[Mux.scala 31:69:@14068.4]
  wire  _T_1643; // @[package.scala 96:25:@14197.4 package.scala 96:25:@14198.4]
  wire [31:0] _T_1647; // @[Mux.scala 31:69:@14207.4]
  wire  _T_1640; // @[package.scala 96:25:@14189.4 package.scala 96:25:@14190.4]
  wire [31:0] _T_1648; // @[Mux.scala 31:69:@14208.4]
  wire  _T_1637; // @[package.scala 96:25:@14181.4 package.scala 96:25:@14182.4]
  wire [31:0] _T_1649; // @[Mux.scala 31:69:@14209.4]
  wire  _T_1634; // @[package.scala 96:25:@14173.4 package.scala 96:25:@14174.4]
  wire [31:0] _T_1650; // @[Mux.scala 31:69:@14210.4]
  wire  _T_1631; // @[package.scala 96:25:@14165.4 package.scala 96:25:@14166.4]
  wire [31:0] _T_1651; // @[Mux.scala 31:69:@14211.4]
  wire  _T_1628; // @[package.scala 96:25:@14157.4 package.scala 96:25:@14158.4]
  wire [31:0] _T_1652; // @[Mux.scala 31:69:@14212.4]
  wire  _T_1625; // @[package.scala 96:25:@14149.4 package.scala 96:25:@14150.4]
  wire [31:0] _T_1653; // @[Mux.scala 31:69:@14213.4]
  wire  _T_1622; // @[package.scala 96:25:@14141.4 package.scala 96:25:@14142.4]
  wire [31:0] _T_1654; // @[Mux.scala 31:69:@14214.4]
  wire  _T_1619; // @[package.scala 96:25:@14133.4 package.scala 96:25:@14134.4]
  wire [31:0] _T_1655; // @[Mux.scala 31:69:@14215.4]
  wire  _T_1616; // @[package.scala 96:25:@14125.4 package.scala 96:25:@14126.4]
  wire [31:0] _T_1656; // @[Mux.scala 31:69:@14216.4]
  wire  _T_1613; // @[package.scala 96:25:@14117.4 package.scala 96:25:@14118.4]
  wire  _T_1750; // @[package.scala 96:25:@14341.4 package.scala 96:25:@14342.4]
  wire [31:0] _T_1754; // @[Mux.scala 31:69:@14351.4]
  wire  _T_1747; // @[package.scala 96:25:@14333.4 package.scala 96:25:@14334.4]
  wire [31:0] _T_1755; // @[Mux.scala 31:69:@14352.4]
  wire  _T_1744; // @[package.scala 96:25:@14325.4 package.scala 96:25:@14326.4]
  wire [31:0] _T_1756; // @[Mux.scala 31:69:@14353.4]
  wire  _T_1741; // @[package.scala 96:25:@14317.4 package.scala 96:25:@14318.4]
  wire [31:0] _T_1757; // @[Mux.scala 31:69:@14354.4]
  wire  _T_1738; // @[package.scala 96:25:@14309.4 package.scala 96:25:@14310.4]
  wire [31:0] _T_1758; // @[Mux.scala 31:69:@14355.4]
  wire  _T_1735; // @[package.scala 96:25:@14301.4 package.scala 96:25:@14302.4]
  wire [31:0] _T_1759; // @[Mux.scala 31:69:@14356.4]
  wire  _T_1732; // @[package.scala 96:25:@14293.4 package.scala 96:25:@14294.4]
  wire [31:0] _T_1760; // @[Mux.scala 31:69:@14357.4]
  wire  _T_1729; // @[package.scala 96:25:@14285.4 package.scala 96:25:@14286.4]
  wire [31:0] _T_1761; // @[Mux.scala 31:69:@14358.4]
  wire  _T_1726; // @[package.scala 96:25:@14277.4 package.scala 96:25:@14278.4]
  wire [31:0] _T_1762; // @[Mux.scala 31:69:@14359.4]
  wire  _T_1723; // @[package.scala 96:25:@14269.4 package.scala 96:25:@14270.4]
  wire [31:0] _T_1763; // @[Mux.scala 31:69:@14360.4]
  wire  _T_1720; // @[package.scala 96:25:@14261.4 package.scala 96:25:@14262.4]
  wire  _T_1857; // @[package.scala 96:25:@14485.4 package.scala 96:25:@14486.4]
  wire [31:0] _T_1861; // @[Mux.scala 31:69:@14495.4]
  wire  _T_1854; // @[package.scala 96:25:@14477.4 package.scala 96:25:@14478.4]
  wire [31:0] _T_1862; // @[Mux.scala 31:69:@14496.4]
  wire  _T_1851; // @[package.scala 96:25:@14469.4 package.scala 96:25:@14470.4]
  wire [31:0] _T_1863; // @[Mux.scala 31:69:@14497.4]
  wire  _T_1848; // @[package.scala 96:25:@14461.4 package.scala 96:25:@14462.4]
  wire [31:0] _T_1864; // @[Mux.scala 31:69:@14498.4]
  wire  _T_1845; // @[package.scala 96:25:@14453.4 package.scala 96:25:@14454.4]
  wire [31:0] _T_1865; // @[Mux.scala 31:69:@14499.4]
  wire  _T_1842; // @[package.scala 96:25:@14445.4 package.scala 96:25:@14446.4]
  wire [31:0] _T_1866; // @[Mux.scala 31:69:@14500.4]
  wire  _T_1839; // @[package.scala 96:25:@14437.4 package.scala 96:25:@14438.4]
  wire [31:0] _T_1867; // @[Mux.scala 31:69:@14501.4]
  wire  _T_1836; // @[package.scala 96:25:@14429.4 package.scala 96:25:@14430.4]
  wire [31:0] _T_1868; // @[Mux.scala 31:69:@14502.4]
  wire  _T_1833; // @[package.scala 96:25:@14421.4 package.scala 96:25:@14422.4]
  wire [31:0] _T_1869; // @[Mux.scala 31:69:@14503.4]
  wire  _T_1830; // @[package.scala 96:25:@14413.4 package.scala 96:25:@14414.4]
  wire [31:0] _T_1870; // @[Mux.scala 31:69:@14504.4]
  wire  _T_1827; // @[package.scala 96:25:@14405.4 package.scala 96:25:@14406.4]
  wire  _T_1964; // @[package.scala 96:25:@14629.4 package.scala 96:25:@14630.4]
  wire [31:0] _T_1968; // @[Mux.scala 31:69:@14639.4]
  wire  _T_1961; // @[package.scala 96:25:@14621.4 package.scala 96:25:@14622.4]
  wire [31:0] _T_1969; // @[Mux.scala 31:69:@14640.4]
  wire  _T_1958; // @[package.scala 96:25:@14613.4 package.scala 96:25:@14614.4]
  wire [31:0] _T_1970; // @[Mux.scala 31:69:@14641.4]
  wire  _T_1955; // @[package.scala 96:25:@14605.4 package.scala 96:25:@14606.4]
  wire [31:0] _T_1971; // @[Mux.scala 31:69:@14642.4]
  wire  _T_1952; // @[package.scala 96:25:@14597.4 package.scala 96:25:@14598.4]
  wire [31:0] _T_1972; // @[Mux.scala 31:69:@14643.4]
  wire  _T_1949; // @[package.scala 96:25:@14589.4 package.scala 96:25:@14590.4]
  wire [31:0] _T_1973; // @[Mux.scala 31:69:@14644.4]
  wire  _T_1946; // @[package.scala 96:25:@14581.4 package.scala 96:25:@14582.4]
  wire [31:0] _T_1974; // @[Mux.scala 31:69:@14645.4]
  wire  _T_1943; // @[package.scala 96:25:@14573.4 package.scala 96:25:@14574.4]
  wire [31:0] _T_1975; // @[Mux.scala 31:69:@14646.4]
  wire  _T_1940; // @[package.scala 96:25:@14565.4 package.scala 96:25:@14566.4]
  wire [31:0] _T_1976; // @[Mux.scala 31:69:@14647.4]
  wire  _T_1937; // @[package.scala 96:25:@14557.4 package.scala 96:25:@14558.4]
  wire [31:0] _T_1977; // @[Mux.scala 31:69:@14648.4]
  wire  _T_1934; // @[package.scala 96:25:@14549.4 package.scala 96:25:@14550.4]
  wire  _T_2071; // @[package.scala 96:25:@14773.4 package.scala 96:25:@14774.4]
  wire [31:0] _T_2075; // @[Mux.scala 31:69:@14783.4]
  wire  _T_2068; // @[package.scala 96:25:@14765.4 package.scala 96:25:@14766.4]
  wire [31:0] _T_2076; // @[Mux.scala 31:69:@14784.4]
  wire  _T_2065; // @[package.scala 96:25:@14757.4 package.scala 96:25:@14758.4]
  wire [31:0] _T_2077; // @[Mux.scala 31:69:@14785.4]
  wire  _T_2062; // @[package.scala 96:25:@14749.4 package.scala 96:25:@14750.4]
  wire [31:0] _T_2078; // @[Mux.scala 31:69:@14786.4]
  wire  _T_2059; // @[package.scala 96:25:@14741.4 package.scala 96:25:@14742.4]
  wire [31:0] _T_2079; // @[Mux.scala 31:69:@14787.4]
  wire  _T_2056; // @[package.scala 96:25:@14733.4 package.scala 96:25:@14734.4]
  wire [31:0] _T_2080; // @[Mux.scala 31:69:@14788.4]
  wire  _T_2053; // @[package.scala 96:25:@14725.4 package.scala 96:25:@14726.4]
  wire [31:0] _T_2081; // @[Mux.scala 31:69:@14789.4]
  wire  _T_2050; // @[package.scala 96:25:@14717.4 package.scala 96:25:@14718.4]
  wire [31:0] _T_2082; // @[Mux.scala 31:69:@14790.4]
  wire  _T_2047; // @[package.scala 96:25:@14709.4 package.scala 96:25:@14710.4]
  wire [31:0] _T_2083; // @[Mux.scala 31:69:@14791.4]
  wire  _T_2044; // @[package.scala 96:25:@14701.4 package.scala 96:25:@14702.4]
  wire [31:0] _T_2084; // @[Mux.scala 31:69:@14792.4]
  wire  _T_2041; // @[package.scala 96:25:@14693.4 package.scala 96:25:@14694.4]
  wire  _T_2178; // @[package.scala 96:25:@14917.4 package.scala 96:25:@14918.4]
  wire [31:0] _T_2182; // @[Mux.scala 31:69:@14927.4]
  wire  _T_2175; // @[package.scala 96:25:@14909.4 package.scala 96:25:@14910.4]
  wire [31:0] _T_2183; // @[Mux.scala 31:69:@14928.4]
  wire  _T_2172; // @[package.scala 96:25:@14901.4 package.scala 96:25:@14902.4]
  wire [31:0] _T_2184; // @[Mux.scala 31:69:@14929.4]
  wire  _T_2169; // @[package.scala 96:25:@14893.4 package.scala 96:25:@14894.4]
  wire [31:0] _T_2185; // @[Mux.scala 31:69:@14930.4]
  wire  _T_2166; // @[package.scala 96:25:@14885.4 package.scala 96:25:@14886.4]
  wire [31:0] _T_2186; // @[Mux.scala 31:69:@14931.4]
  wire  _T_2163; // @[package.scala 96:25:@14877.4 package.scala 96:25:@14878.4]
  wire [31:0] _T_2187; // @[Mux.scala 31:69:@14932.4]
  wire  _T_2160; // @[package.scala 96:25:@14869.4 package.scala 96:25:@14870.4]
  wire [31:0] _T_2188; // @[Mux.scala 31:69:@14933.4]
  wire  _T_2157; // @[package.scala 96:25:@14861.4 package.scala 96:25:@14862.4]
  wire [31:0] _T_2189; // @[Mux.scala 31:69:@14934.4]
  wire  _T_2154; // @[package.scala 96:25:@14853.4 package.scala 96:25:@14854.4]
  wire [31:0] _T_2190; // @[Mux.scala 31:69:@14935.4]
  wire  _T_2151; // @[package.scala 96:25:@14845.4 package.scala 96:25:@14846.4]
  wire [31:0] _T_2191; // @[Mux.scala 31:69:@14936.4]
  wire  _T_2148; // @[package.scala 96:25:@14837.4 package.scala 96:25:@14838.4]
  wire  _T_2285; // @[package.scala 96:25:@15061.4 package.scala 96:25:@15062.4]
  wire [31:0] _T_2289; // @[Mux.scala 31:69:@15071.4]
  wire  _T_2282; // @[package.scala 96:25:@15053.4 package.scala 96:25:@15054.4]
  wire [31:0] _T_2290; // @[Mux.scala 31:69:@15072.4]
  wire  _T_2279; // @[package.scala 96:25:@15045.4 package.scala 96:25:@15046.4]
  wire [31:0] _T_2291; // @[Mux.scala 31:69:@15073.4]
  wire  _T_2276; // @[package.scala 96:25:@15037.4 package.scala 96:25:@15038.4]
  wire [31:0] _T_2292; // @[Mux.scala 31:69:@15074.4]
  wire  _T_2273; // @[package.scala 96:25:@15029.4 package.scala 96:25:@15030.4]
  wire [31:0] _T_2293; // @[Mux.scala 31:69:@15075.4]
  wire  _T_2270; // @[package.scala 96:25:@15021.4 package.scala 96:25:@15022.4]
  wire [31:0] _T_2294; // @[Mux.scala 31:69:@15076.4]
  wire  _T_2267; // @[package.scala 96:25:@15013.4 package.scala 96:25:@15014.4]
  wire [31:0] _T_2295; // @[Mux.scala 31:69:@15077.4]
  wire  _T_2264; // @[package.scala 96:25:@15005.4 package.scala 96:25:@15006.4]
  wire [31:0] _T_2296; // @[Mux.scala 31:69:@15078.4]
  wire  _T_2261; // @[package.scala 96:25:@14997.4 package.scala 96:25:@14998.4]
  wire [31:0] _T_2297; // @[Mux.scala 31:69:@15079.4]
  wire  _T_2258; // @[package.scala 96:25:@14989.4 package.scala 96:25:@14990.4]
  wire [31:0] _T_2298; // @[Mux.scala 31:69:@15080.4]
  wire  _T_2255; // @[package.scala 96:25:@14981.4 package.scala 96:25:@14982.4]
  wire  _T_2392; // @[package.scala 96:25:@15205.4 package.scala 96:25:@15206.4]
  wire [31:0] _T_2396; // @[Mux.scala 31:69:@15215.4]
  wire  _T_2389; // @[package.scala 96:25:@15197.4 package.scala 96:25:@15198.4]
  wire [31:0] _T_2397; // @[Mux.scala 31:69:@15216.4]
  wire  _T_2386; // @[package.scala 96:25:@15189.4 package.scala 96:25:@15190.4]
  wire [31:0] _T_2398; // @[Mux.scala 31:69:@15217.4]
  wire  _T_2383; // @[package.scala 96:25:@15181.4 package.scala 96:25:@15182.4]
  wire [31:0] _T_2399; // @[Mux.scala 31:69:@15218.4]
  wire  _T_2380; // @[package.scala 96:25:@15173.4 package.scala 96:25:@15174.4]
  wire [31:0] _T_2400; // @[Mux.scala 31:69:@15219.4]
  wire  _T_2377; // @[package.scala 96:25:@15165.4 package.scala 96:25:@15166.4]
  wire [31:0] _T_2401; // @[Mux.scala 31:69:@15220.4]
  wire  _T_2374; // @[package.scala 96:25:@15157.4 package.scala 96:25:@15158.4]
  wire [31:0] _T_2402; // @[Mux.scala 31:69:@15221.4]
  wire  _T_2371; // @[package.scala 96:25:@15149.4 package.scala 96:25:@15150.4]
  wire [31:0] _T_2403; // @[Mux.scala 31:69:@15222.4]
  wire  _T_2368; // @[package.scala 96:25:@15141.4 package.scala 96:25:@15142.4]
  wire [31:0] _T_2404; // @[Mux.scala 31:69:@15223.4]
  wire  _T_2365; // @[package.scala 96:25:@15133.4 package.scala 96:25:@15134.4]
  wire [31:0] _T_2405; // @[Mux.scala 31:69:@15224.4]
  wire  _T_2362; // @[package.scala 96:25:@15125.4 package.scala 96:25:@15126.4]
  wire  _T_2499; // @[package.scala 96:25:@15349.4 package.scala 96:25:@15350.4]
  wire [31:0] _T_2503; // @[Mux.scala 31:69:@15359.4]
  wire  _T_2496; // @[package.scala 96:25:@15341.4 package.scala 96:25:@15342.4]
  wire [31:0] _T_2504; // @[Mux.scala 31:69:@15360.4]
  wire  _T_2493; // @[package.scala 96:25:@15333.4 package.scala 96:25:@15334.4]
  wire [31:0] _T_2505; // @[Mux.scala 31:69:@15361.4]
  wire  _T_2490; // @[package.scala 96:25:@15325.4 package.scala 96:25:@15326.4]
  wire [31:0] _T_2506; // @[Mux.scala 31:69:@15362.4]
  wire  _T_2487; // @[package.scala 96:25:@15317.4 package.scala 96:25:@15318.4]
  wire [31:0] _T_2507; // @[Mux.scala 31:69:@15363.4]
  wire  _T_2484; // @[package.scala 96:25:@15309.4 package.scala 96:25:@15310.4]
  wire [31:0] _T_2508; // @[Mux.scala 31:69:@15364.4]
  wire  _T_2481; // @[package.scala 96:25:@15301.4 package.scala 96:25:@15302.4]
  wire [31:0] _T_2509; // @[Mux.scala 31:69:@15365.4]
  wire  _T_2478; // @[package.scala 96:25:@15293.4 package.scala 96:25:@15294.4]
  wire [31:0] _T_2510; // @[Mux.scala 31:69:@15366.4]
  wire  _T_2475; // @[package.scala 96:25:@15285.4 package.scala 96:25:@15286.4]
  wire [31:0] _T_2511; // @[Mux.scala 31:69:@15367.4]
  wire  _T_2472; // @[package.scala 96:25:@15277.4 package.scala 96:25:@15278.4]
  wire [31:0] _T_2512; // @[Mux.scala 31:69:@15368.4]
  wire  _T_2469; // @[package.scala 96:25:@15269.4 package.scala 96:25:@15270.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12671.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12687.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12703.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12719.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12735.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12751.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12767.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12783.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12799.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12815.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12831.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12847.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@13043.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@13132.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@13221.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13310.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13399.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13488.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13577.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13666.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13755.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13844.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13933.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@14022.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@14112.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@14120.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@14128.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@14136.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@14144.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@14152.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@14160.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@14168.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@14176.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@14184.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@14192.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14200.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14256.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14264.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14272.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14280.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14288.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14296.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14304.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14312.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14320.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14328.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14336.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14344.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14400.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14408.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14416.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14424.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14432.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14440.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14448.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14456.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14464.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14472.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14480.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14488.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14544.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14552.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14560.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14568.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14576.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14584.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14592.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14600.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14608.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14616.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14624.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14632.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14688.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14696.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14704.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14712.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14720.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14728.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14736.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14744.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14752.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14760.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14768.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14776.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14832.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14840.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14848.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14856.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14864.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14872.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14880.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@14888.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@14896.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@14904.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@14912.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@14920.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@14976.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@14984.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@14992.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@15000.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@15008.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@15016.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@15024.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@15032.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@15040.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@15048.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@15056.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@15064.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@15120.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@15128.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@15136.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@15144.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@15152.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@15160.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@15168.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@15176.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@15184.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@15192.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15200.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15208.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@15264.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@15272.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@15280.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@15288.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@15296.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@15304.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@15312.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@15320.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@15328.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@15336.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@15344.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@15352.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  assign _T_316 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12863.4]
  assign _T_318 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@12864.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 82:228:@12865.4]
  assign _T_320 = io_wPort_0_en_0 & _T_319; // @[MemPrimitives.scala 83:102:@12866.4]
  assign _T_322 = {_T_320,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12868.4]
  assign _T_329 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@12876.4]
  assign _T_330 = _T_316 & _T_329; // @[MemPrimitives.scala 82:228:@12877.4]
  assign _T_331 = io_wPort_0_en_0 & _T_330; // @[MemPrimitives.scala 83:102:@12878.4]
  assign _T_333 = {_T_331,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12880.4]
  assign _T_340 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@12888.4]
  assign _T_341 = _T_316 & _T_340; // @[MemPrimitives.scala 82:228:@12889.4]
  assign _T_342 = io_wPort_0_en_0 & _T_341; // @[MemPrimitives.scala 83:102:@12890.4]
  assign _T_344 = {_T_342,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12892.4]
  assign _T_349 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12899.4]
  assign _T_352 = _T_349 & _T_318; // @[MemPrimitives.scala 82:228:@12901.4]
  assign _T_353 = io_wPort_0_en_0 & _T_352; // @[MemPrimitives.scala 83:102:@12902.4]
  assign _T_355 = {_T_353,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12904.4]
  assign _T_363 = _T_349 & _T_329; // @[MemPrimitives.scala 82:228:@12913.4]
  assign _T_364 = io_wPort_0_en_0 & _T_363; // @[MemPrimitives.scala 83:102:@12914.4]
  assign _T_366 = {_T_364,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12916.4]
  assign _T_374 = _T_349 & _T_340; // @[MemPrimitives.scala 82:228:@12925.4]
  assign _T_375 = io_wPort_0_en_0 & _T_374; // @[MemPrimitives.scala 83:102:@12926.4]
  assign _T_377 = {_T_375,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12928.4]
  assign _T_382 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12935.4]
  assign _T_385 = _T_382 & _T_318; // @[MemPrimitives.scala 82:228:@12937.4]
  assign _T_386 = io_wPort_0_en_0 & _T_385; // @[MemPrimitives.scala 83:102:@12938.4]
  assign _T_388 = {_T_386,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12940.4]
  assign _T_396 = _T_382 & _T_329; // @[MemPrimitives.scala 82:228:@12949.4]
  assign _T_397 = io_wPort_0_en_0 & _T_396; // @[MemPrimitives.scala 83:102:@12950.4]
  assign _T_399 = {_T_397,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12952.4]
  assign _T_407 = _T_382 & _T_340; // @[MemPrimitives.scala 82:228:@12961.4]
  assign _T_408 = io_wPort_0_en_0 & _T_407; // @[MemPrimitives.scala 83:102:@12962.4]
  assign _T_410 = {_T_408,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12964.4]
  assign _T_415 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12971.4]
  assign _T_418 = _T_415 & _T_318; // @[MemPrimitives.scala 82:228:@12973.4]
  assign _T_419 = io_wPort_0_en_0 & _T_418; // @[MemPrimitives.scala 83:102:@12974.4]
  assign _T_421 = {_T_419,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12976.4]
  assign _T_429 = _T_415 & _T_329; // @[MemPrimitives.scala 82:228:@12985.4]
  assign _T_430 = io_wPort_0_en_0 & _T_429; // @[MemPrimitives.scala 83:102:@12986.4]
  assign _T_432 = {_T_430,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12988.4]
  assign _T_440 = _T_415 & _T_340; // @[MemPrimitives.scala 82:228:@12997.4]
  assign _T_441 = io_wPort_0_en_0 & _T_440; // @[MemPrimitives.scala 83:102:@12998.4]
  assign _T_443 = {_T_441,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13000.4]
  assign _T_448 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13007.4]
  assign _T_450 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13008.4]
  assign _T_451 = _T_448 & _T_450; // @[MemPrimitives.scala 110:228:@13009.4]
  assign _T_454 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13011.4]
  assign _T_456 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13012.4]
  assign _T_457 = _T_454 & _T_456; // @[MemPrimitives.scala 110:228:@13013.4]
  assign _T_460 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13015.4]
  assign _T_462 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13016.4]
  assign _T_463 = _T_460 & _T_462; // @[MemPrimitives.scala 110:228:@13017.4]
  assign _T_466 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13019.4]
  assign _T_468 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13020.4]
  assign _T_469 = _T_466 & _T_468; // @[MemPrimitives.scala 110:228:@13021.4]
  assign _T_472 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13023.4]
  assign _T_474 = io_rPort_4_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13024.4]
  assign _T_475 = _T_472 & _T_474; // @[MemPrimitives.scala 110:228:@13025.4]
  assign _T_478 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13027.4]
  assign _T_480 = io_rPort_5_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13028.4]
  assign _T_481 = _T_478 & _T_480; // @[MemPrimitives.scala 110:228:@13029.4]
  assign _T_484 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13031.4]
  assign _T_486 = io_rPort_6_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13032.4]
  assign _T_487 = _T_484 & _T_486; // @[MemPrimitives.scala 110:228:@13033.4]
  assign _T_490 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13035.4]
  assign _T_492 = io_rPort_7_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13036.4]
  assign _T_493 = _T_490 & _T_492; // @[MemPrimitives.scala 110:228:@13037.4]
  assign _T_496 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13039.4]
  assign _T_498 = io_rPort_8_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13040.4]
  assign _T_499 = _T_496 & _T_498; // @[MemPrimitives.scala 110:228:@13041.4]
  assign _T_501 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@13055.4]
  assign _T_502 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@13056.4]
  assign _T_503 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@13057.4]
  assign _T_504 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@13058.4]
  assign _T_505 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@13059.4]
  assign _T_506 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@13060.4]
  assign _T_507 = StickySelects_io_outs_6; // @[MemPrimitives.scala 126:35:@13061.4]
  assign _T_508 = StickySelects_io_outs_7; // @[MemPrimitives.scala 126:35:@13062.4]
  assign _T_509 = StickySelects_io_outs_8; // @[MemPrimitives.scala 126:35:@13063.4]
  assign _T_511 = {_T_501,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13065.4]
  assign _T_513 = {_T_502,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13067.4]
  assign _T_515 = {_T_503,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13069.4]
  assign _T_517 = {_T_504,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13071.4]
  assign _T_519 = {_T_505,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13073.4]
  assign _T_521 = {_T_506,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13075.4]
  assign _T_523 = {_T_507,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13077.4]
  assign _T_525 = {_T_508,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13079.4]
  assign _T_527 = {_T_509,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13081.4]
  assign _T_528 = _T_508 ? _T_525 : _T_527; // @[Mux.scala 31:69:@13082.4]
  assign _T_529 = _T_507 ? _T_523 : _T_528; // @[Mux.scala 31:69:@13083.4]
  assign _T_530 = _T_506 ? _T_521 : _T_529; // @[Mux.scala 31:69:@13084.4]
  assign _T_531 = _T_505 ? _T_519 : _T_530; // @[Mux.scala 31:69:@13085.4]
  assign _T_532 = _T_504 ? _T_517 : _T_531; // @[Mux.scala 31:69:@13086.4]
  assign _T_533 = _T_503 ? _T_515 : _T_532; // @[Mux.scala 31:69:@13087.4]
  assign _T_534 = _T_502 ? _T_513 : _T_533; // @[Mux.scala 31:69:@13088.4]
  assign _T_535 = _T_501 ? _T_511 : _T_534; // @[Mux.scala 31:69:@13089.4]
  assign _T_542 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13097.4]
  assign _T_543 = _T_448 & _T_542; // @[MemPrimitives.scala 110:228:@13098.4]
  assign _T_548 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13101.4]
  assign _T_549 = _T_454 & _T_548; // @[MemPrimitives.scala 110:228:@13102.4]
  assign _T_554 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13105.4]
  assign _T_555 = _T_460 & _T_554; // @[MemPrimitives.scala 110:228:@13106.4]
  assign _T_560 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13109.4]
  assign _T_561 = _T_466 & _T_560; // @[MemPrimitives.scala 110:228:@13110.4]
  assign _T_566 = io_rPort_4_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13113.4]
  assign _T_567 = _T_472 & _T_566; // @[MemPrimitives.scala 110:228:@13114.4]
  assign _T_572 = io_rPort_5_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13117.4]
  assign _T_573 = _T_478 & _T_572; // @[MemPrimitives.scala 110:228:@13118.4]
  assign _T_578 = io_rPort_6_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13121.4]
  assign _T_579 = _T_484 & _T_578; // @[MemPrimitives.scala 110:228:@13122.4]
  assign _T_584 = io_rPort_7_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13125.4]
  assign _T_585 = _T_490 & _T_584; // @[MemPrimitives.scala 110:228:@13126.4]
  assign _T_590 = io_rPort_8_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13129.4]
  assign _T_591 = _T_496 & _T_590; // @[MemPrimitives.scala 110:228:@13130.4]
  assign _T_593 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@13144.4]
  assign _T_594 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@13145.4]
  assign _T_595 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@13146.4]
  assign _T_596 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@13147.4]
  assign _T_597 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@13148.4]
  assign _T_598 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@13149.4]
  assign _T_599 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 126:35:@13150.4]
  assign _T_600 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 126:35:@13151.4]
  assign _T_601 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 126:35:@13152.4]
  assign _T_603 = {_T_593,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13154.4]
  assign _T_605 = {_T_594,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13156.4]
  assign _T_607 = {_T_595,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13158.4]
  assign _T_609 = {_T_596,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13160.4]
  assign _T_611 = {_T_597,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13162.4]
  assign _T_613 = {_T_598,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13164.4]
  assign _T_615 = {_T_599,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13166.4]
  assign _T_617 = {_T_600,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13168.4]
  assign _T_619 = {_T_601,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13170.4]
  assign _T_620 = _T_600 ? _T_617 : _T_619; // @[Mux.scala 31:69:@13171.4]
  assign _T_621 = _T_599 ? _T_615 : _T_620; // @[Mux.scala 31:69:@13172.4]
  assign _T_622 = _T_598 ? _T_613 : _T_621; // @[Mux.scala 31:69:@13173.4]
  assign _T_623 = _T_597 ? _T_611 : _T_622; // @[Mux.scala 31:69:@13174.4]
  assign _T_624 = _T_596 ? _T_609 : _T_623; // @[Mux.scala 31:69:@13175.4]
  assign _T_625 = _T_595 ? _T_607 : _T_624; // @[Mux.scala 31:69:@13176.4]
  assign _T_626 = _T_594 ? _T_605 : _T_625; // @[Mux.scala 31:69:@13177.4]
  assign _T_627 = _T_593 ? _T_603 : _T_626; // @[Mux.scala 31:69:@13178.4]
  assign _T_634 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13186.4]
  assign _T_635 = _T_448 & _T_634; // @[MemPrimitives.scala 110:228:@13187.4]
  assign _T_640 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13190.4]
  assign _T_641 = _T_454 & _T_640; // @[MemPrimitives.scala 110:228:@13191.4]
  assign _T_646 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13194.4]
  assign _T_647 = _T_460 & _T_646; // @[MemPrimitives.scala 110:228:@13195.4]
  assign _T_652 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13198.4]
  assign _T_653 = _T_466 & _T_652; // @[MemPrimitives.scala 110:228:@13199.4]
  assign _T_658 = io_rPort_4_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13202.4]
  assign _T_659 = _T_472 & _T_658; // @[MemPrimitives.scala 110:228:@13203.4]
  assign _T_664 = io_rPort_5_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13206.4]
  assign _T_665 = _T_478 & _T_664; // @[MemPrimitives.scala 110:228:@13207.4]
  assign _T_670 = io_rPort_6_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13210.4]
  assign _T_671 = _T_484 & _T_670; // @[MemPrimitives.scala 110:228:@13211.4]
  assign _T_676 = io_rPort_7_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13214.4]
  assign _T_677 = _T_490 & _T_676; // @[MemPrimitives.scala 110:228:@13215.4]
  assign _T_682 = io_rPort_8_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13218.4]
  assign _T_683 = _T_496 & _T_682; // @[MemPrimitives.scala 110:228:@13219.4]
  assign _T_685 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@13233.4]
  assign _T_686 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@13234.4]
  assign _T_687 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@13235.4]
  assign _T_688 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@13236.4]
  assign _T_689 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@13237.4]
  assign _T_690 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@13238.4]
  assign _T_691 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 126:35:@13239.4]
  assign _T_692 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 126:35:@13240.4]
  assign _T_693 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 126:35:@13241.4]
  assign _T_695 = {_T_685,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13243.4]
  assign _T_697 = {_T_686,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13245.4]
  assign _T_699 = {_T_687,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13247.4]
  assign _T_701 = {_T_688,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13249.4]
  assign _T_703 = {_T_689,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13251.4]
  assign _T_705 = {_T_690,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13253.4]
  assign _T_707 = {_T_691,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13255.4]
  assign _T_709 = {_T_692,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13257.4]
  assign _T_711 = {_T_693,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13259.4]
  assign _T_712 = _T_692 ? _T_709 : _T_711; // @[Mux.scala 31:69:@13260.4]
  assign _T_713 = _T_691 ? _T_707 : _T_712; // @[Mux.scala 31:69:@13261.4]
  assign _T_714 = _T_690 ? _T_705 : _T_713; // @[Mux.scala 31:69:@13262.4]
  assign _T_715 = _T_689 ? _T_703 : _T_714; // @[Mux.scala 31:69:@13263.4]
  assign _T_716 = _T_688 ? _T_701 : _T_715; // @[Mux.scala 31:69:@13264.4]
  assign _T_717 = _T_687 ? _T_699 : _T_716; // @[Mux.scala 31:69:@13265.4]
  assign _T_718 = _T_686 ? _T_697 : _T_717; // @[Mux.scala 31:69:@13266.4]
  assign _T_719 = _T_685 ? _T_695 : _T_718; // @[Mux.scala 31:69:@13267.4]
  assign _T_724 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13274.4]
  assign _T_727 = _T_724 & _T_450; // @[MemPrimitives.scala 110:228:@13276.4]
  assign _T_730 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13278.4]
  assign _T_733 = _T_730 & _T_456; // @[MemPrimitives.scala 110:228:@13280.4]
  assign _T_736 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13282.4]
  assign _T_739 = _T_736 & _T_462; // @[MemPrimitives.scala 110:228:@13284.4]
  assign _T_742 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13286.4]
  assign _T_745 = _T_742 & _T_468; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_748 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13290.4]
  assign _T_751 = _T_748 & _T_474; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_754 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13294.4]
  assign _T_757 = _T_754 & _T_480; // @[MemPrimitives.scala 110:228:@13296.4]
  assign _T_760 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13298.4]
  assign _T_763 = _T_760 & _T_486; // @[MemPrimitives.scala 110:228:@13300.4]
  assign _T_766 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13302.4]
  assign _T_769 = _T_766 & _T_492; // @[MemPrimitives.scala 110:228:@13304.4]
  assign _T_772 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13306.4]
  assign _T_775 = _T_772 & _T_498; // @[MemPrimitives.scala 110:228:@13308.4]
  assign _T_777 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13322.4]
  assign _T_778 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13323.4]
  assign _T_779 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13324.4]
  assign _T_780 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13325.4]
  assign _T_781 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13326.4]
  assign _T_782 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13327.4]
  assign _T_783 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 126:35:@13328.4]
  assign _T_784 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 126:35:@13329.4]
  assign _T_785 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 126:35:@13330.4]
  assign _T_787 = {_T_777,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13332.4]
  assign _T_789 = {_T_778,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13334.4]
  assign _T_791 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13336.4]
  assign _T_793 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13338.4]
  assign _T_795 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13340.4]
  assign _T_797 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13342.4]
  assign _T_799 = {_T_783,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13344.4]
  assign _T_801 = {_T_784,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13346.4]
  assign _T_803 = {_T_785,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13348.4]
  assign _T_804 = _T_784 ? _T_801 : _T_803; // @[Mux.scala 31:69:@13349.4]
  assign _T_805 = _T_783 ? _T_799 : _T_804; // @[Mux.scala 31:69:@13350.4]
  assign _T_806 = _T_782 ? _T_797 : _T_805; // @[Mux.scala 31:69:@13351.4]
  assign _T_807 = _T_781 ? _T_795 : _T_806; // @[Mux.scala 31:69:@13352.4]
  assign _T_808 = _T_780 ? _T_793 : _T_807; // @[Mux.scala 31:69:@13353.4]
  assign _T_809 = _T_779 ? _T_791 : _T_808; // @[Mux.scala 31:69:@13354.4]
  assign _T_810 = _T_778 ? _T_789 : _T_809; // @[Mux.scala 31:69:@13355.4]
  assign _T_811 = _T_777 ? _T_787 : _T_810; // @[Mux.scala 31:69:@13356.4]
  assign _T_819 = _T_724 & _T_542; // @[MemPrimitives.scala 110:228:@13365.4]
  assign _T_825 = _T_730 & _T_548; // @[MemPrimitives.scala 110:228:@13369.4]
  assign _T_831 = _T_736 & _T_554; // @[MemPrimitives.scala 110:228:@13373.4]
  assign _T_837 = _T_742 & _T_560; // @[MemPrimitives.scala 110:228:@13377.4]
  assign _T_843 = _T_748 & _T_566; // @[MemPrimitives.scala 110:228:@13381.4]
  assign _T_849 = _T_754 & _T_572; // @[MemPrimitives.scala 110:228:@13385.4]
  assign _T_855 = _T_760 & _T_578; // @[MemPrimitives.scala 110:228:@13389.4]
  assign _T_861 = _T_766 & _T_584; // @[MemPrimitives.scala 110:228:@13393.4]
  assign _T_867 = _T_772 & _T_590; // @[MemPrimitives.scala 110:228:@13397.4]
  assign _T_869 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13411.4]
  assign _T_870 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13412.4]
  assign _T_871 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13413.4]
  assign _T_872 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13414.4]
  assign _T_873 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13415.4]
  assign _T_874 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13416.4]
  assign _T_875 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 126:35:@13417.4]
  assign _T_876 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 126:35:@13418.4]
  assign _T_877 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 126:35:@13419.4]
  assign _T_879 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13421.4]
  assign _T_881 = {_T_870,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13423.4]
  assign _T_883 = {_T_871,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13425.4]
  assign _T_885 = {_T_872,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13427.4]
  assign _T_887 = {_T_873,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13429.4]
  assign _T_889 = {_T_874,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13431.4]
  assign _T_891 = {_T_875,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13433.4]
  assign _T_893 = {_T_876,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13435.4]
  assign _T_895 = {_T_877,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13437.4]
  assign _T_896 = _T_876 ? _T_893 : _T_895; // @[Mux.scala 31:69:@13438.4]
  assign _T_897 = _T_875 ? _T_891 : _T_896; // @[Mux.scala 31:69:@13439.4]
  assign _T_898 = _T_874 ? _T_889 : _T_897; // @[Mux.scala 31:69:@13440.4]
  assign _T_899 = _T_873 ? _T_887 : _T_898; // @[Mux.scala 31:69:@13441.4]
  assign _T_900 = _T_872 ? _T_885 : _T_899; // @[Mux.scala 31:69:@13442.4]
  assign _T_901 = _T_871 ? _T_883 : _T_900; // @[Mux.scala 31:69:@13443.4]
  assign _T_902 = _T_870 ? _T_881 : _T_901; // @[Mux.scala 31:69:@13444.4]
  assign _T_903 = _T_869 ? _T_879 : _T_902; // @[Mux.scala 31:69:@13445.4]
  assign _T_911 = _T_724 & _T_634; // @[MemPrimitives.scala 110:228:@13454.4]
  assign _T_917 = _T_730 & _T_640; // @[MemPrimitives.scala 110:228:@13458.4]
  assign _T_923 = _T_736 & _T_646; // @[MemPrimitives.scala 110:228:@13462.4]
  assign _T_929 = _T_742 & _T_652; // @[MemPrimitives.scala 110:228:@13466.4]
  assign _T_935 = _T_748 & _T_658; // @[MemPrimitives.scala 110:228:@13470.4]
  assign _T_941 = _T_754 & _T_664; // @[MemPrimitives.scala 110:228:@13474.4]
  assign _T_947 = _T_760 & _T_670; // @[MemPrimitives.scala 110:228:@13478.4]
  assign _T_953 = _T_766 & _T_676; // @[MemPrimitives.scala 110:228:@13482.4]
  assign _T_959 = _T_772 & _T_682; // @[MemPrimitives.scala 110:228:@13486.4]
  assign _T_961 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13500.4]
  assign _T_962 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13501.4]
  assign _T_963 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13502.4]
  assign _T_964 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13503.4]
  assign _T_965 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13504.4]
  assign _T_966 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13505.4]
  assign _T_967 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 126:35:@13506.4]
  assign _T_968 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 126:35:@13507.4]
  assign _T_969 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 126:35:@13508.4]
  assign _T_971 = {_T_961,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13510.4]
  assign _T_973 = {_T_962,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13512.4]
  assign _T_975 = {_T_963,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13514.4]
  assign _T_977 = {_T_964,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13516.4]
  assign _T_979 = {_T_965,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13518.4]
  assign _T_981 = {_T_966,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13520.4]
  assign _T_983 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13522.4]
  assign _T_985 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13524.4]
  assign _T_987 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13526.4]
  assign _T_988 = _T_968 ? _T_985 : _T_987; // @[Mux.scala 31:69:@13527.4]
  assign _T_989 = _T_967 ? _T_983 : _T_988; // @[Mux.scala 31:69:@13528.4]
  assign _T_990 = _T_966 ? _T_981 : _T_989; // @[Mux.scala 31:69:@13529.4]
  assign _T_991 = _T_965 ? _T_979 : _T_990; // @[Mux.scala 31:69:@13530.4]
  assign _T_992 = _T_964 ? _T_977 : _T_991; // @[Mux.scala 31:69:@13531.4]
  assign _T_993 = _T_963 ? _T_975 : _T_992; // @[Mux.scala 31:69:@13532.4]
  assign _T_994 = _T_962 ? _T_973 : _T_993; // @[Mux.scala 31:69:@13533.4]
  assign _T_995 = _T_961 ? _T_971 : _T_994; // @[Mux.scala 31:69:@13534.4]
  assign _T_1000 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13541.4]
  assign _T_1003 = _T_1000 & _T_450; // @[MemPrimitives.scala 110:228:@13543.4]
  assign _T_1006 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13545.4]
  assign _T_1009 = _T_1006 & _T_456; // @[MemPrimitives.scala 110:228:@13547.4]
  assign _T_1012 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13549.4]
  assign _T_1015 = _T_1012 & _T_462; // @[MemPrimitives.scala 110:228:@13551.4]
  assign _T_1018 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13553.4]
  assign _T_1021 = _T_1018 & _T_468; // @[MemPrimitives.scala 110:228:@13555.4]
  assign _T_1024 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13557.4]
  assign _T_1027 = _T_1024 & _T_474; // @[MemPrimitives.scala 110:228:@13559.4]
  assign _T_1030 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13561.4]
  assign _T_1033 = _T_1030 & _T_480; // @[MemPrimitives.scala 110:228:@13563.4]
  assign _T_1036 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13565.4]
  assign _T_1039 = _T_1036 & _T_486; // @[MemPrimitives.scala 110:228:@13567.4]
  assign _T_1042 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13569.4]
  assign _T_1045 = _T_1042 & _T_492; // @[MemPrimitives.scala 110:228:@13571.4]
  assign _T_1048 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13573.4]
  assign _T_1051 = _T_1048 & _T_498; // @[MemPrimitives.scala 110:228:@13575.4]
  assign _T_1053 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13589.4]
  assign _T_1054 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13590.4]
  assign _T_1055 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13591.4]
  assign _T_1056 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13592.4]
  assign _T_1057 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13593.4]
  assign _T_1058 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13594.4]
  assign _T_1059 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 126:35:@13595.4]
  assign _T_1060 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 126:35:@13596.4]
  assign _T_1061 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 126:35:@13597.4]
  assign _T_1063 = {_T_1053,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13599.4]
  assign _T_1065 = {_T_1054,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13601.4]
  assign _T_1067 = {_T_1055,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13603.4]
  assign _T_1069 = {_T_1056,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13605.4]
  assign _T_1071 = {_T_1057,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13607.4]
  assign _T_1073 = {_T_1058,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13609.4]
  assign _T_1075 = {_T_1059,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13611.4]
  assign _T_1077 = {_T_1060,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13613.4]
  assign _T_1079 = {_T_1061,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13615.4]
  assign _T_1080 = _T_1060 ? _T_1077 : _T_1079; // @[Mux.scala 31:69:@13616.4]
  assign _T_1081 = _T_1059 ? _T_1075 : _T_1080; // @[Mux.scala 31:69:@13617.4]
  assign _T_1082 = _T_1058 ? _T_1073 : _T_1081; // @[Mux.scala 31:69:@13618.4]
  assign _T_1083 = _T_1057 ? _T_1071 : _T_1082; // @[Mux.scala 31:69:@13619.4]
  assign _T_1084 = _T_1056 ? _T_1069 : _T_1083; // @[Mux.scala 31:69:@13620.4]
  assign _T_1085 = _T_1055 ? _T_1067 : _T_1084; // @[Mux.scala 31:69:@13621.4]
  assign _T_1086 = _T_1054 ? _T_1065 : _T_1085; // @[Mux.scala 31:69:@13622.4]
  assign _T_1087 = _T_1053 ? _T_1063 : _T_1086; // @[Mux.scala 31:69:@13623.4]
  assign _T_1095 = _T_1000 & _T_542; // @[MemPrimitives.scala 110:228:@13632.4]
  assign _T_1101 = _T_1006 & _T_548; // @[MemPrimitives.scala 110:228:@13636.4]
  assign _T_1107 = _T_1012 & _T_554; // @[MemPrimitives.scala 110:228:@13640.4]
  assign _T_1113 = _T_1018 & _T_560; // @[MemPrimitives.scala 110:228:@13644.4]
  assign _T_1119 = _T_1024 & _T_566; // @[MemPrimitives.scala 110:228:@13648.4]
  assign _T_1125 = _T_1030 & _T_572; // @[MemPrimitives.scala 110:228:@13652.4]
  assign _T_1131 = _T_1036 & _T_578; // @[MemPrimitives.scala 110:228:@13656.4]
  assign _T_1137 = _T_1042 & _T_584; // @[MemPrimitives.scala 110:228:@13660.4]
  assign _T_1143 = _T_1048 & _T_590; // @[MemPrimitives.scala 110:228:@13664.4]
  assign _T_1145 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13678.4]
  assign _T_1146 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13679.4]
  assign _T_1147 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13680.4]
  assign _T_1148 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13681.4]
  assign _T_1149 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13682.4]
  assign _T_1150 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13683.4]
  assign _T_1151 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 126:35:@13684.4]
  assign _T_1152 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 126:35:@13685.4]
  assign _T_1153 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 126:35:@13686.4]
  assign _T_1155 = {_T_1145,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13688.4]
  assign _T_1157 = {_T_1146,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13690.4]
  assign _T_1159 = {_T_1147,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13692.4]
  assign _T_1161 = {_T_1148,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13694.4]
  assign _T_1163 = {_T_1149,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13696.4]
  assign _T_1165 = {_T_1150,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13698.4]
  assign _T_1167 = {_T_1151,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13700.4]
  assign _T_1169 = {_T_1152,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13702.4]
  assign _T_1171 = {_T_1153,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13704.4]
  assign _T_1172 = _T_1152 ? _T_1169 : _T_1171; // @[Mux.scala 31:69:@13705.4]
  assign _T_1173 = _T_1151 ? _T_1167 : _T_1172; // @[Mux.scala 31:69:@13706.4]
  assign _T_1174 = _T_1150 ? _T_1165 : _T_1173; // @[Mux.scala 31:69:@13707.4]
  assign _T_1175 = _T_1149 ? _T_1163 : _T_1174; // @[Mux.scala 31:69:@13708.4]
  assign _T_1176 = _T_1148 ? _T_1161 : _T_1175; // @[Mux.scala 31:69:@13709.4]
  assign _T_1177 = _T_1147 ? _T_1159 : _T_1176; // @[Mux.scala 31:69:@13710.4]
  assign _T_1178 = _T_1146 ? _T_1157 : _T_1177; // @[Mux.scala 31:69:@13711.4]
  assign _T_1179 = _T_1145 ? _T_1155 : _T_1178; // @[Mux.scala 31:69:@13712.4]
  assign _T_1187 = _T_1000 & _T_634; // @[MemPrimitives.scala 110:228:@13721.4]
  assign _T_1193 = _T_1006 & _T_640; // @[MemPrimitives.scala 110:228:@13725.4]
  assign _T_1199 = _T_1012 & _T_646; // @[MemPrimitives.scala 110:228:@13729.4]
  assign _T_1205 = _T_1018 & _T_652; // @[MemPrimitives.scala 110:228:@13733.4]
  assign _T_1211 = _T_1024 & _T_658; // @[MemPrimitives.scala 110:228:@13737.4]
  assign _T_1217 = _T_1030 & _T_664; // @[MemPrimitives.scala 110:228:@13741.4]
  assign _T_1223 = _T_1036 & _T_670; // @[MemPrimitives.scala 110:228:@13745.4]
  assign _T_1229 = _T_1042 & _T_676; // @[MemPrimitives.scala 110:228:@13749.4]
  assign _T_1235 = _T_1048 & _T_682; // @[MemPrimitives.scala 110:228:@13753.4]
  assign _T_1237 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13767.4]
  assign _T_1238 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13768.4]
  assign _T_1239 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13769.4]
  assign _T_1240 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13770.4]
  assign _T_1241 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13771.4]
  assign _T_1242 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13772.4]
  assign _T_1243 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 126:35:@13773.4]
  assign _T_1244 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 126:35:@13774.4]
  assign _T_1245 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 126:35:@13775.4]
  assign _T_1247 = {_T_1237,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13777.4]
  assign _T_1249 = {_T_1238,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13779.4]
  assign _T_1251 = {_T_1239,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13781.4]
  assign _T_1253 = {_T_1240,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13783.4]
  assign _T_1255 = {_T_1241,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13785.4]
  assign _T_1257 = {_T_1242,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13787.4]
  assign _T_1259 = {_T_1243,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13789.4]
  assign _T_1261 = {_T_1244,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13791.4]
  assign _T_1263 = {_T_1245,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13793.4]
  assign _T_1264 = _T_1244 ? _T_1261 : _T_1263; // @[Mux.scala 31:69:@13794.4]
  assign _T_1265 = _T_1243 ? _T_1259 : _T_1264; // @[Mux.scala 31:69:@13795.4]
  assign _T_1266 = _T_1242 ? _T_1257 : _T_1265; // @[Mux.scala 31:69:@13796.4]
  assign _T_1267 = _T_1241 ? _T_1255 : _T_1266; // @[Mux.scala 31:69:@13797.4]
  assign _T_1268 = _T_1240 ? _T_1253 : _T_1267; // @[Mux.scala 31:69:@13798.4]
  assign _T_1269 = _T_1239 ? _T_1251 : _T_1268; // @[Mux.scala 31:69:@13799.4]
  assign _T_1270 = _T_1238 ? _T_1249 : _T_1269; // @[Mux.scala 31:69:@13800.4]
  assign _T_1271 = _T_1237 ? _T_1247 : _T_1270; // @[Mux.scala 31:69:@13801.4]
  assign _T_1276 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13808.4]
  assign _T_1279 = _T_1276 & _T_450; // @[MemPrimitives.scala 110:228:@13810.4]
  assign _T_1282 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13812.4]
  assign _T_1285 = _T_1282 & _T_456; // @[MemPrimitives.scala 110:228:@13814.4]
  assign _T_1288 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13816.4]
  assign _T_1291 = _T_1288 & _T_462; // @[MemPrimitives.scala 110:228:@13818.4]
  assign _T_1294 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13820.4]
  assign _T_1297 = _T_1294 & _T_468; // @[MemPrimitives.scala 110:228:@13822.4]
  assign _T_1300 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13824.4]
  assign _T_1303 = _T_1300 & _T_474; // @[MemPrimitives.scala 110:228:@13826.4]
  assign _T_1306 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13828.4]
  assign _T_1309 = _T_1306 & _T_480; // @[MemPrimitives.scala 110:228:@13830.4]
  assign _T_1312 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13832.4]
  assign _T_1315 = _T_1312 & _T_486; // @[MemPrimitives.scala 110:228:@13834.4]
  assign _T_1318 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13836.4]
  assign _T_1321 = _T_1318 & _T_492; // @[MemPrimitives.scala 110:228:@13838.4]
  assign _T_1324 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13840.4]
  assign _T_1327 = _T_1324 & _T_498; // @[MemPrimitives.scala 110:228:@13842.4]
  assign _T_1329 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13856.4]
  assign _T_1330 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13857.4]
  assign _T_1331 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13858.4]
  assign _T_1332 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13859.4]
  assign _T_1333 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13860.4]
  assign _T_1334 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13861.4]
  assign _T_1335 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 126:35:@13862.4]
  assign _T_1336 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 126:35:@13863.4]
  assign _T_1337 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 126:35:@13864.4]
  assign _T_1339 = {_T_1329,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13866.4]
  assign _T_1341 = {_T_1330,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13868.4]
  assign _T_1343 = {_T_1331,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13870.4]
  assign _T_1345 = {_T_1332,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13872.4]
  assign _T_1347 = {_T_1333,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13874.4]
  assign _T_1349 = {_T_1334,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13876.4]
  assign _T_1351 = {_T_1335,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13878.4]
  assign _T_1353 = {_T_1336,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13880.4]
  assign _T_1355 = {_T_1337,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13882.4]
  assign _T_1356 = _T_1336 ? _T_1353 : _T_1355; // @[Mux.scala 31:69:@13883.4]
  assign _T_1357 = _T_1335 ? _T_1351 : _T_1356; // @[Mux.scala 31:69:@13884.4]
  assign _T_1358 = _T_1334 ? _T_1349 : _T_1357; // @[Mux.scala 31:69:@13885.4]
  assign _T_1359 = _T_1333 ? _T_1347 : _T_1358; // @[Mux.scala 31:69:@13886.4]
  assign _T_1360 = _T_1332 ? _T_1345 : _T_1359; // @[Mux.scala 31:69:@13887.4]
  assign _T_1361 = _T_1331 ? _T_1343 : _T_1360; // @[Mux.scala 31:69:@13888.4]
  assign _T_1362 = _T_1330 ? _T_1341 : _T_1361; // @[Mux.scala 31:69:@13889.4]
  assign _T_1363 = _T_1329 ? _T_1339 : _T_1362; // @[Mux.scala 31:69:@13890.4]
  assign _T_1371 = _T_1276 & _T_542; // @[MemPrimitives.scala 110:228:@13899.4]
  assign _T_1377 = _T_1282 & _T_548; // @[MemPrimitives.scala 110:228:@13903.4]
  assign _T_1383 = _T_1288 & _T_554; // @[MemPrimitives.scala 110:228:@13907.4]
  assign _T_1389 = _T_1294 & _T_560; // @[MemPrimitives.scala 110:228:@13911.4]
  assign _T_1395 = _T_1300 & _T_566; // @[MemPrimitives.scala 110:228:@13915.4]
  assign _T_1401 = _T_1306 & _T_572; // @[MemPrimitives.scala 110:228:@13919.4]
  assign _T_1407 = _T_1312 & _T_578; // @[MemPrimitives.scala 110:228:@13923.4]
  assign _T_1413 = _T_1318 & _T_584; // @[MemPrimitives.scala 110:228:@13927.4]
  assign _T_1419 = _T_1324 & _T_590; // @[MemPrimitives.scala 110:228:@13931.4]
  assign _T_1421 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13945.4]
  assign _T_1422 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13946.4]
  assign _T_1423 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13947.4]
  assign _T_1424 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13948.4]
  assign _T_1425 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13949.4]
  assign _T_1426 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13950.4]
  assign _T_1427 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 126:35:@13951.4]
  assign _T_1428 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 126:35:@13952.4]
  assign _T_1429 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 126:35:@13953.4]
  assign _T_1431 = {_T_1421,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13955.4]
  assign _T_1433 = {_T_1422,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13957.4]
  assign _T_1435 = {_T_1423,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13959.4]
  assign _T_1437 = {_T_1424,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13961.4]
  assign _T_1439 = {_T_1425,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13963.4]
  assign _T_1441 = {_T_1426,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13965.4]
  assign _T_1443 = {_T_1427,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13967.4]
  assign _T_1445 = {_T_1428,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13969.4]
  assign _T_1447 = {_T_1429,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13971.4]
  assign _T_1448 = _T_1428 ? _T_1445 : _T_1447; // @[Mux.scala 31:69:@13972.4]
  assign _T_1449 = _T_1427 ? _T_1443 : _T_1448; // @[Mux.scala 31:69:@13973.4]
  assign _T_1450 = _T_1426 ? _T_1441 : _T_1449; // @[Mux.scala 31:69:@13974.4]
  assign _T_1451 = _T_1425 ? _T_1439 : _T_1450; // @[Mux.scala 31:69:@13975.4]
  assign _T_1452 = _T_1424 ? _T_1437 : _T_1451; // @[Mux.scala 31:69:@13976.4]
  assign _T_1453 = _T_1423 ? _T_1435 : _T_1452; // @[Mux.scala 31:69:@13977.4]
  assign _T_1454 = _T_1422 ? _T_1433 : _T_1453; // @[Mux.scala 31:69:@13978.4]
  assign _T_1455 = _T_1421 ? _T_1431 : _T_1454; // @[Mux.scala 31:69:@13979.4]
  assign _T_1463 = _T_1276 & _T_634; // @[MemPrimitives.scala 110:228:@13988.4]
  assign _T_1469 = _T_1282 & _T_640; // @[MemPrimitives.scala 110:228:@13992.4]
  assign _T_1475 = _T_1288 & _T_646; // @[MemPrimitives.scala 110:228:@13996.4]
  assign _T_1481 = _T_1294 & _T_652; // @[MemPrimitives.scala 110:228:@14000.4]
  assign _T_1487 = _T_1300 & _T_658; // @[MemPrimitives.scala 110:228:@14004.4]
  assign _T_1493 = _T_1306 & _T_664; // @[MemPrimitives.scala 110:228:@14008.4]
  assign _T_1499 = _T_1312 & _T_670; // @[MemPrimitives.scala 110:228:@14012.4]
  assign _T_1505 = _T_1318 & _T_676; // @[MemPrimitives.scala 110:228:@14016.4]
  assign _T_1511 = _T_1324 & _T_682; // @[MemPrimitives.scala 110:228:@14020.4]
  assign _T_1513 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@14034.4]
  assign _T_1514 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@14035.4]
  assign _T_1515 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@14036.4]
  assign _T_1516 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@14037.4]
  assign _T_1517 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@14038.4]
  assign _T_1518 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@14039.4]
  assign _T_1519 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 126:35:@14040.4]
  assign _T_1520 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 126:35:@14041.4]
  assign _T_1521 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 126:35:@14042.4]
  assign _T_1523 = {_T_1513,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14044.4]
  assign _T_1525 = {_T_1514,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14046.4]
  assign _T_1527 = {_T_1515,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14048.4]
  assign _T_1529 = {_T_1516,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14050.4]
  assign _T_1531 = {_T_1517,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14052.4]
  assign _T_1533 = {_T_1518,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14054.4]
  assign _T_1535 = {_T_1519,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14056.4]
  assign _T_1537 = {_T_1520,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14058.4]
  assign _T_1539 = {_T_1521,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14060.4]
  assign _T_1540 = _T_1520 ? _T_1537 : _T_1539; // @[Mux.scala 31:69:@14061.4]
  assign _T_1541 = _T_1519 ? _T_1535 : _T_1540; // @[Mux.scala 31:69:@14062.4]
  assign _T_1542 = _T_1518 ? _T_1533 : _T_1541; // @[Mux.scala 31:69:@14063.4]
  assign _T_1543 = _T_1517 ? _T_1531 : _T_1542; // @[Mux.scala 31:69:@14064.4]
  assign _T_1544 = _T_1516 ? _T_1529 : _T_1543; // @[Mux.scala 31:69:@14065.4]
  assign _T_1545 = _T_1515 ? _T_1527 : _T_1544; // @[Mux.scala 31:69:@14066.4]
  assign _T_1546 = _T_1514 ? _T_1525 : _T_1545; // @[Mux.scala 31:69:@14067.4]
  assign _T_1547 = _T_1513 ? _T_1523 : _T_1546; // @[Mux.scala 31:69:@14068.4]
  assign _T_1643 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14197.4 package.scala 96:25:@14198.4]
  assign _T_1647 = _T_1643 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14207.4]
  assign _T_1640 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14189.4 package.scala 96:25:@14190.4]
  assign _T_1648 = _T_1640 ? Mem1D_9_io_output : _T_1647; // @[Mux.scala 31:69:@14208.4]
  assign _T_1637 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14181.4 package.scala 96:25:@14182.4]
  assign _T_1649 = _T_1637 ? Mem1D_8_io_output : _T_1648; // @[Mux.scala 31:69:@14209.4]
  assign _T_1634 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@14173.4 package.scala 96:25:@14174.4]
  assign _T_1650 = _T_1634 ? Mem1D_7_io_output : _T_1649; // @[Mux.scala 31:69:@14210.4]
  assign _T_1631 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14165.4 package.scala 96:25:@14166.4]
  assign _T_1651 = _T_1631 ? Mem1D_6_io_output : _T_1650; // @[Mux.scala 31:69:@14211.4]
  assign _T_1628 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14157.4 package.scala 96:25:@14158.4]
  assign _T_1652 = _T_1628 ? Mem1D_5_io_output : _T_1651; // @[Mux.scala 31:69:@14212.4]
  assign _T_1625 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14149.4 package.scala 96:25:@14150.4]
  assign _T_1653 = _T_1625 ? Mem1D_4_io_output : _T_1652; // @[Mux.scala 31:69:@14213.4]
  assign _T_1622 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14141.4 package.scala 96:25:@14142.4]
  assign _T_1654 = _T_1622 ? Mem1D_3_io_output : _T_1653; // @[Mux.scala 31:69:@14214.4]
  assign _T_1619 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14133.4 package.scala 96:25:@14134.4]
  assign _T_1655 = _T_1619 ? Mem1D_2_io_output : _T_1654; // @[Mux.scala 31:69:@14215.4]
  assign _T_1616 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14125.4 package.scala 96:25:@14126.4]
  assign _T_1656 = _T_1616 ? Mem1D_1_io_output : _T_1655; // @[Mux.scala 31:69:@14216.4]
  assign _T_1613 = RetimeWrapper_io_out; // @[package.scala 96:25:@14117.4 package.scala 96:25:@14118.4]
  assign _T_1750 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14341.4 package.scala 96:25:@14342.4]
  assign _T_1754 = _T_1750 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14351.4]
  assign _T_1747 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14333.4 package.scala 96:25:@14334.4]
  assign _T_1755 = _T_1747 ? Mem1D_9_io_output : _T_1754; // @[Mux.scala 31:69:@14352.4]
  assign _T_1744 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14325.4 package.scala 96:25:@14326.4]
  assign _T_1756 = _T_1744 ? Mem1D_8_io_output : _T_1755; // @[Mux.scala 31:69:@14353.4]
  assign _T_1741 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14317.4 package.scala 96:25:@14318.4]
  assign _T_1757 = _T_1741 ? Mem1D_7_io_output : _T_1756; // @[Mux.scala 31:69:@14354.4]
  assign _T_1738 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14309.4 package.scala 96:25:@14310.4]
  assign _T_1758 = _T_1738 ? Mem1D_6_io_output : _T_1757; // @[Mux.scala 31:69:@14355.4]
  assign _T_1735 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14301.4 package.scala 96:25:@14302.4]
  assign _T_1759 = _T_1735 ? Mem1D_5_io_output : _T_1758; // @[Mux.scala 31:69:@14356.4]
  assign _T_1732 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14293.4 package.scala 96:25:@14294.4]
  assign _T_1760 = _T_1732 ? Mem1D_4_io_output : _T_1759; // @[Mux.scala 31:69:@14357.4]
  assign _T_1729 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@14285.4 package.scala 96:25:@14286.4]
  assign _T_1761 = _T_1729 ? Mem1D_3_io_output : _T_1760; // @[Mux.scala 31:69:@14358.4]
  assign _T_1726 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14277.4 package.scala 96:25:@14278.4]
  assign _T_1762 = _T_1726 ? Mem1D_2_io_output : _T_1761; // @[Mux.scala 31:69:@14359.4]
  assign _T_1723 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14269.4 package.scala 96:25:@14270.4]
  assign _T_1763 = _T_1723 ? Mem1D_1_io_output : _T_1762; // @[Mux.scala 31:69:@14360.4]
  assign _T_1720 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14261.4 package.scala 96:25:@14262.4]
  assign _T_1857 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14485.4 package.scala 96:25:@14486.4]
  assign _T_1861 = _T_1857 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14495.4]
  assign _T_1854 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14477.4 package.scala 96:25:@14478.4]
  assign _T_1862 = _T_1854 ? Mem1D_9_io_output : _T_1861; // @[Mux.scala 31:69:@14496.4]
  assign _T_1851 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14469.4 package.scala 96:25:@14470.4]
  assign _T_1863 = _T_1851 ? Mem1D_8_io_output : _T_1862; // @[Mux.scala 31:69:@14497.4]
  assign _T_1848 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@14461.4 package.scala 96:25:@14462.4]
  assign _T_1864 = _T_1848 ? Mem1D_7_io_output : _T_1863; // @[Mux.scala 31:69:@14498.4]
  assign _T_1845 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14453.4 package.scala 96:25:@14454.4]
  assign _T_1865 = _T_1845 ? Mem1D_6_io_output : _T_1864; // @[Mux.scala 31:69:@14499.4]
  assign _T_1842 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14445.4 package.scala 96:25:@14446.4]
  assign _T_1866 = _T_1842 ? Mem1D_5_io_output : _T_1865; // @[Mux.scala 31:69:@14500.4]
  assign _T_1839 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14437.4 package.scala 96:25:@14438.4]
  assign _T_1867 = _T_1839 ? Mem1D_4_io_output : _T_1866; // @[Mux.scala 31:69:@14501.4]
  assign _T_1836 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14429.4 package.scala 96:25:@14430.4]
  assign _T_1868 = _T_1836 ? Mem1D_3_io_output : _T_1867; // @[Mux.scala 31:69:@14502.4]
  assign _T_1833 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14421.4 package.scala 96:25:@14422.4]
  assign _T_1869 = _T_1833 ? Mem1D_2_io_output : _T_1868; // @[Mux.scala 31:69:@14503.4]
  assign _T_1830 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14413.4 package.scala 96:25:@14414.4]
  assign _T_1870 = _T_1830 ? Mem1D_1_io_output : _T_1869; // @[Mux.scala 31:69:@14504.4]
  assign _T_1827 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14405.4 package.scala 96:25:@14406.4]
  assign _T_1964 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14629.4 package.scala 96:25:@14630.4]
  assign _T_1968 = _T_1964 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14639.4]
  assign _T_1961 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14621.4 package.scala 96:25:@14622.4]
  assign _T_1969 = _T_1961 ? Mem1D_9_io_output : _T_1968; // @[Mux.scala 31:69:@14640.4]
  assign _T_1958 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14613.4 package.scala 96:25:@14614.4]
  assign _T_1970 = _T_1958 ? Mem1D_8_io_output : _T_1969; // @[Mux.scala 31:69:@14641.4]
  assign _T_1955 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14605.4 package.scala 96:25:@14606.4]
  assign _T_1971 = _T_1955 ? Mem1D_7_io_output : _T_1970; // @[Mux.scala 31:69:@14642.4]
  assign _T_1952 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14597.4 package.scala 96:25:@14598.4]
  assign _T_1972 = _T_1952 ? Mem1D_6_io_output : _T_1971; // @[Mux.scala 31:69:@14643.4]
  assign _T_1949 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14589.4 package.scala 96:25:@14590.4]
  assign _T_1973 = _T_1949 ? Mem1D_5_io_output : _T_1972; // @[Mux.scala 31:69:@14644.4]
  assign _T_1946 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14581.4 package.scala 96:25:@14582.4]
  assign _T_1974 = _T_1946 ? Mem1D_4_io_output : _T_1973; // @[Mux.scala 31:69:@14645.4]
  assign _T_1943 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@14573.4 package.scala 96:25:@14574.4]
  assign _T_1975 = _T_1943 ? Mem1D_3_io_output : _T_1974; // @[Mux.scala 31:69:@14646.4]
  assign _T_1940 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14565.4 package.scala 96:25:@14566.4]
  assign _T_1976 = _T_1940 ? Mem1D_2_io_output : _T_1975; // @[Mux.scala 31:69:@14647.4]
  assign _T_1937 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14557.4 package.scala 96:25:@14558.4]
  assign _T_1977 = _T_1937 ? Mem1D_1_io_output : _T_1976; // @[Mux.scala 31:69:@14648.4]
  assign _T_1934 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14549.4 package.scala 96:25:@14550.4]
  assign _T_2071 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14773.4 package.scala 96:25:@14774.4]
  assign _T_2075 = _T_2071 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14783.4]
  assign _T_2068 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14765.4 package.scala 96:25:@14766.4]
  assign _T_2076 = _T_2068 ? Mem1D_9_io_output : _T_2075; // @[Mux.scala 31:69:@14784.4]
  assign _T_2065 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14757.4 package.scala 96:25:@14758.4]
  assign _T_2077 = _T_2065 ? Mem1D_8_io_output : _T_2076; // @[Mux.scala 31:69:@14785.4]
  assign _T_2062 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@14749.4 package.scala 96:25:@14750.4]
  assign _T_2078 = _T_2062 ? Mem1D_7_io_output : _T_2077; // @[Mux.scala 31:69:@14786.4]
  assign _T_2059 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14741.4 package.scala 96:25:@14742.4]
  assign _T_2079 = _T_2059 ? Mem1D_6_io_output : _T_2078; // @[Mux.scala 31:69:@14787.4]
  assign _T_2056 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14733.4 package.scala 96:25:@14734.4]
  assign _T_2080 = _T_2056 ? Mem1D_5_io_output : _T_2079; // @[Mux.scala 31:69:@14788.4]
  assign _T_2053 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14725.4 package.scala 96:25:@14726.4]
  assign _T_2081 = _T_2053 ? Mem1D_4_io_output : _T_2080; // @[Mux.scala 31:69:@14789.4]
  assign _T_2050 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14717.4 package.scala 96:25:@14718.4]
  assign _T_2082 = _T_2050 ? Mem1D_3_io_output : _T_2081; // @[Mux.scala 31:69:@14790.4]
  assign _T_2047 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14709.4 package.scala 96:25:@14710.4]
  assign _T_2083 = _T_2047 ? Mem1D_2_io_output : _T_2082; // @[Mux.scala 31:69:@14791.4]
  assign _T_2044 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14701.4 package.scala 96:25:@14702.4]
  assign _T_2084 = _T_2044 ? Mem1D_1_io_output : _T_2083; // @[Mux.scala 31:69:@14792.4]
  assign _T_2041 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14693.4 package.scala 96:25:@14694.4]
  assign _T_2178 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14917.4 package.scala 96:25:@14918.4]
  assign _T_2182 = _T_2178 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14927.4]
  assign _T_2175 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14909.4 package.scala 96:25:@14910.4]
  assign _T_2183 = _T_2175 ? Mem1D_9_io_output : _T_2182; // @[Mux.scala 31:69:@14928.4]
  assign _T_2172 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14901.4 package.scala 96:25:@14902.4]
  assign _T_2184 = _T_2172 ? Mem1D_8_io_output : _T_2183; // @[Mux.scala 31:69:@14929.4]
  assign _T_2169 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14893.4 package.scala 96:25:@14894.4]
  assign _T_2185 = _T_2169 ? Mem1D_7_io_output : _T_2184; // @[Mux.scala 31:69:@14930.4]
  assign _T_2166 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14885.4 package.scala 96:25:@14886.4]
  assign _T_2186 = _T_2166 ? Mem1D_6_io_output : _T_2185; // @[Mux.scala 31:69:@14931.4]
  assign _T_2163 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14877.4 package.scala 96:25:@14878.4]
  assign _T_2187 = _T_2163 ? Mem1D_5_io_output : _T_2186; // @[Mux.scala 31:69:@14932.4]
  assign _T_2160 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14869.4 package.scala 96:25:@14870.4]
  assign _T_2188 = _T_2160 ? Mem1D_4_io_output : _T_2187; // @[Mux.scala 31:69:@14933.4]
  assign _T_2157 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@14861.4 package.scala 96:25:@14862.4]
  assign _T_2189 = _T_2157 ? Mem1D_3_io_output : _T_2188; // @[Mux.scala 31:69:@14934.4]
  assign _T_2154 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14853.4 package.scala 96:25:@14854.4]
  assign _T_2190 = _T_2154 ? Mem1D_2_io_output : _T_2189; // @[Mux.scala 31:69:@14935.4]
  assign _T_2151 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14845.4 package.scala 96:25:@14846.4]
  assign _T_2191 = _T_2151 ? Mem1D_1_io_output : _T_2190; // @[Mux.scala 31:69:@14936.4]
  assign _T_2148 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14837.4 package.scala 96:25:@14838.4]
  assign _T_2285 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@15061.4 package.scala 96:25:@15062.4]
  assign _T_2289 = _T_2285 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15071.4]
  assign _T_2282 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@15053.4 package.scala 96:25:@15054.4]
  assign _T_2290 = _T_2282 ? Mem1D_9_io_output : _T_2289; // @[Mux.scala 31:69:@15072.4]
  assign _T_2279 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@15045.4 package.scala 96:25:@15046.4]
  assign _T_2291 = _T_2279 ? Mem1D_8_io_output : _T_2290; // @[Mux.scala 31:69:@15073.4]
  assign _T_2276 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@15037.4 package.scala 96:25:@15038.4]
  assign _T_2292 = _T_2276 ? Mem1D_7_io_output : _T_2291; // @[Mux.scala 31:69:@15074.4]
  assign _T_2273 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@15029.4 package.scala 96:25:@15030.4]
  assign _T_2293 = _T_2273 ? Mem1D_6_io_output : _T_2292; // @[Mux.scala 31:69:@15075.4]
  assign _T_2270 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@15021.4 package.scala 96:25:@15022.4]
  assign _T_2294 = _T_2270 ? Mem1D_5_io_output : _T_2293; // @[Mux.scala 31:69:@15076.4]
  assign _T_2267 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@15013.4 package.scala 96:25:@15014.4]
  assign _T_2295 = _T_2267 ? Mem1D_4_io_output : _T_2294; // @[Mux.scala 31:69:@15077.4]
  assign _T_2264 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@15005.4 package.scala 96:25:@15006.4]
  assign _T_2296 = _T_2264 ? Mem1D_3_io_output : _T_2295; // @[Mux.scala 31:69:@15078.4]
  assign _T_2261 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14997.4 package.scala 96:25:@14998.4]
  assign _T_2297 = _T_2261 ? Mem1D_2_io_output : _T_2296; // @[Mux.scala 31:69:@15079.4]
  assign _T_2258 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14989.4 package.scala 96:25:@14990.4]
  assign _T_2298 = _T_2258 ? Mem1D_1_io_output : _T_2297; // @[Mux.scala 31:69:@15080.4]
  assign _T_2255 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14981.4 package.scala 96:25:@14982.4]
  assign _T_2392 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15205.4 package.scala 96:25:@15206.4]
  assign _T_2396 = _T_2392 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15215.4]
  assign _T_2389 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15197.4 package.scala 96:25:@15198.4]
  assign _T_2397 = _T_2389 ? Mem1D_9_io_output : _T_2396; // @[Mux.scala 31:69:@15216.4]
  assign _T_2386 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@15189.4 package.scala 96:25:@15190.4]
  assign _T_2398 = _T_2386 ? Mem1D_8_io_output : _T_2397; // @[Mux.scala 31:69:@15217.4]
  assign _T_2383 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@15181.4 package.scala 96:25:@15182.4]
  assign _T_2399 = _T_2383 ? Mem1D_7_io_output : _T_2398; // @[Mux.scala 31:69:@15218.4]
  assign _T_2380 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@15173.4 package.scala 96:25:@15174.4]
  assign _T_2400 = _T_2380 ? Mem1D_6_io_output : _T_2399; // @[Mux.scala 31:69:@15219.4]
  assign _T_2377 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@15165.4 package.scala 96:25:@15166.4]
  assign _T_2401 = _T_2377 ? Mem1D_5_io_output : _T_2400; // @[Mux.scala 31:69:@15220.4]
  assign _T_2374 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@15157.4 package.scala 96:25:@15158.4]
  assign _T_2402 = _T_2374 ? Mem1D_4_io_output : _T_2401; // @[Mux.scala 31:69:@15221.4]
  assign _T_2371 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@15149.4 package.scala 96:25:@15150.4]
  assign _T_2403 = _T_2371 ? Mem1D_3_io_output : _T_2402; // @[Mux.scala 31:69:@15222.4]
  assign _T_2368 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@15141.4 package.scala 96:25:@15142.4]
  assign _T_2404 = _T_2368 ? Mem1D_2_io_output : _T_2403; // @[Mux.scala 31:69:@15223.4]
  assign _T_2365 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@15133.4 package.scala 96:25:@15134.4]
  assign _T_2405 = _T_2365 ? Mem1D_1_io_output : _T_2404; // @[Mux.scala 31:69:@15224.4]
  assign _T_2362 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@15125.4 package.scala 96:25:@15126.4]
  assign _T_2499 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@15349.4 package.scala 96:25:@15350.4]
  assign _T_2503 = _T_2499 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15359.4]
  assign _T_2496 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@15341.4 package.scala 96:25:@15342.4]
  assign _T_2504 = _T_2496 ? Mem1D_9_io_output : _T_2503; // @[Mux.scala 31:69:@15360.4]
  assign _T_2493 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@15333.4 package.scala 96:25:@15334.4]
  assign _T_2505 = _T_2493 ? Mem1D_8_io_output : _T_2504; // @[Mux.scala 31:69:@15361.4]
  assign _T_2490 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@15325.4 package.scala 96:25:@15326.4]
  assign _T_2506 = _T_2490 ? Mem1D_7_io_output : _T_2505; // @[Mux.scala 31:69:@15362.4]
  assign _T_2487 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@15317.4 package.scala 96:25:@15318.4]
  assign _T_2507 = _T_2487 ? Mem1D_6_io_output : _T_2506; // @[Mux.scala 31:69:@15363.4]
  assign _T_2484 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@15309.4 package.scala 96:25:@15310.4]
  assign _T_2508 = _T_2484 ? Mem1D_5_io_output : _T_2507; // @[Mux.scala 31:69:@15364.4]
  assign _T_2481 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@15301.4 package.scala 96:25:@15302.4]
  assign _T_2509 = _T_2481 ? Mem1D_4_io_output : _T_2508; // @[Mux.scala 31:69:@15365.4]
  assign _T_2478 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@15293.4 package.scala 96:25:@15294.4]
  assign _T_2510 = _T_2478 ? Mem1D_3_io_output : _T_2509; // @[Mux.scala 31:69:@15366.4]
  assign _T_2475 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@15285.4 package.scala 96:25:@15286.4]
  assign _T_2511 = _T_2475 ? Mem1D_2_io_output : _T_2510; // @[Mux.scala 31:69:@15367.4]
  assign _T_2472 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@15277.4 package.scala 96:25:@15278.4]
  assign _T_2512 = _T_2472 ? Mem1D_1_io_output : _T_2511; // @[Mux.scala 31:69:@15368.4]
  assign _T_2469 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@15269.4 package.scala 96:25:@15270.4]
  assign io_rPort_8_output_0 = _T_2469 ? Mem1D_io_output : _T_2512; // @[MemPrimitives.scala 152:13:@15370.4]
  assign io_rPort_7_output_0 = _T_2362 ? Mem1D_io_output : _T_2405; // @[MemPrimitives.scala 152:13:@15226.4]
  assign io_rPort_6_output_0 = _T_2255 ? Mem1D_io_output : _T_2298; // @[MemPrimitives.scala 152:13:@15082.4]
  assign io_rPort_5_output_0 = _T_2148 ? Mem1D_io_output : _T_2191; // @[MemPrimitives.scala 152:13:@14938.4]
  assign io_rPort_4_output_0 = _T_2041 ? Mem1D_io_output : _T_2084; // @[MemPrimitives.scala 152:13:@14794.4]
  assign io_rPort_3_output_0 = _T_1934 ? Mem1D_io_output : _T_1977; // @[MemPrimitives.scala 152:13:@14650.4]
  assign io_rPort_2_output_0 = _T_1827 ? Mem1D_io_output : _T_1870; // @[MemPrimitives.scala 152:13:@14506.4]
  assign io_rPort_1_output_0 = _T_1720 ? Mem1D_io_output : _T_1763; // @[MemPrimitives.scala 152:13:@14362.4]
  assign io_rPort_0_output_0 = _T_1613 ? Mem1D_io_output : _T_1656; // @[MemPrimitives.scala 152:13:@14218.4]
  assign Mem1D_clock = clock; // @[:@12672.4]
  assign Mem1D_reset = reset; // @[:@12673.4]
  assign Mem1D_io_r_ofs_0 = _T_535[9:0]; // @[MemPrimitives.scala 131:28:@13093.4]
  assign Mem1D_io_r_backpressure = _T_535[10]; // @[MemPrimitives.scala 132:32:@13094.4]
  assign Mem1D_io_w_ofs_0 = _T_322[9:0]; // @[MemPrimitives.scala 94:28:@12872.4]
  assign Mem1D_io_w_data_0 = _T_322[41:10]; // @[MemPrimitives.scala 95:29:@12873.4]
  assign Mem1D_io_w_en_0 = _T_322[42]; // @[MemPrimitives.scala 96:27:@12874.4]
  assign Mem1D_1_clock = clock; // @[:@12688.4]
  assign Mem1D_1_reset = reset; // @[:@12689.4]
  assign Mem1D_1_io_r_ofs_0 = _T_627[9:0]; // @[MemPrimitives.scala 131:28:@13182.4]
  assign Mem1D_1_io_r_backpressure = _T_627[10]; // @[MemPrimitives.scala 132:32:@13183.4]
  assign Mem1D_1_io_w_ofs_0 = _T_333[9:0]; // @[MemPrimitives.scala 94:28:@12884.4]
  assign Mem1D_1_io_w_data_0 = _T_333[41:10]; // @[MemPrimitives.scala 95:29:@12885.4]
  assign Mem1D_1_io_w_en_0 = _T_333[42]; // @[MemPrimitives.scala 96:27:@12886.4]
  assign Mem1D_2_clock = clock; // @[:@12704.4]
  assign Mem1D_2_reset = reset; // @[:@12705.4]
  assign Mem1D_2_io_r_ofs_0 = _T_719[9:0]; // @[MemPrimitives.scala 131:28:@13271.4]
  assign Mem1D_2_io_r_backpressure = _T_719[10]; // @[MemPrimitives.scala 132:32:@13272.4]
  assign Mem1D_2_io_w_ofs_0 = _T_344[9:0]; // @[MemPrimitives.scala 94:28:@12896.4]
  assign Mem1D_2_io_w_data_0 = _T_344[41:10]; // @[MemPrimitives.scala 95:29:@12897.4]
  assign Mem1D_2_io_w_en_0 = _T_344[42]; // @[MemPrimitives.scala 96:27:@12898.4]
  assign Mem1D_3_clock = clock; // @[:@12720.4]
  assign Mem1D_3_reset = reset; // @[:@12721.4]
  assign Mem1D_3_io_r_ofs_0 = _T_811[9:0]; // @[MemPrimitives.scala 131:28:@13360.4]
  assign Mem1D_3_io_r_backpressure = _T_811[10]; // @[MemPrimitives.scala 132:32:@13361.4]
  assign Mem1D_3_io_w_ofs_0 = _T_355[9:0]; // @[MemPrimitives.scala 94:28:@12908.4]
  assign Mem1D_3_io_w_data_0 = _T_355[41:10]; // @[MemPrimitives.scala 95:29:@12909.4]
  assign Mem1D_3_io_w_en_0 = _T_355[42]; // @[MemPrimitives.scala 96:27:@12910.4]
  assign Mem1D_4_clock = clock; // @[:@12736.4]
  assign Mem1D_4_reset = reset; // @[:@12737.4]
  assign Mem1D_4_io_r_ofs_0 = _T_903[9:0]; // @[MemPrimitives.scala 131:28:@13449.4]
  assign Mem1D_4_io_r_backpressure = _T_903[10]; // @[MemPrimitives.scala 132:32:@13450.4]
  assign Mem1D_4_io_w_ofs_0 = _T_366[9:0]; // @[MemPrimitives.scala 94:28:@12920.4]
  assign Mem1D_4_io_w_data_0 = _T_366[41:10]; // @[MemPrimitives.scala 95:29:@12921.4]
  assign Mem1D_4_io_w_en_0 = _T_366[42]; // @[MemPrimitives.scala 96:27:@12922.4]
  assign Mem1D_5_clock = clock; // @[:@12752.4]
  assign Mem1D_5_reset = reset; // @[:@12753.4]
  assign Mem1D_5_io_r_ofs_0 = _T_995[9:0]; // @[MemPrimitives.scala 131:28:@13538.4]
  assign Mem1D_5_io_r_backpressure = _T_995[10]; // @[MemPrimitives.scala 132:32:@13539.4]
  assign Mem1D_5_io_w_ofs_0 = _T_377[9:0]; // @[MemPrimitives.scala 94:28:@12932.4]
  assign Mem1D_5_io_w_data_0 = _T_377[41:10]; // @[MemPrimitives.scala 95:29:@12933.4]
  assign Mem1D_5_io_w_en_0 = _T_377[42]; // @[MemPrimitives.scala 96:27:@12934.4]
  assign Mem1D_6_clock = clock; // @[:@12768.4]
  assign Mem1D_6_reset = reset; // @[:@12769.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1087[9:0]; // @[MemPrimitives.scala 131:28:@13627.4]
  assign Mem1D_6_io_r_backpressure = _T_1087[10]; // @[MemPrimitives.scala 132:32:@13628.4]
  assign Mem1D_6_io_w_ofs_0 = _T_388[9:0]; // @[MemPrimitives.scala 94:28:@12944.4]
  assign Mem1D_6_io_w_data_0 = _T_388[41:10]; // @[MemPrimitives.scala 95:29:@12945.4]
  assign Mem1D_6_io_w_en_0 = _T_388[42]; // @[MemPrimitives.scala 96:27:@12946.4]
  assign Mem1D_7_clock = clock; // @[:@12784.4]
  assign Mem1D_7_reset = reset; // @[:@12785.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1179[9:0]; // @[MemPrimitives.scala 131:28:@13716.4]
  assign Mem1D_7_io_r_backpressure = _T_1179[10]; // @[MemPrimitives.scala 132:32:@13717.4]
  assign Mem1D_7_io_w_ofs_0 = _T_399[9:0]; // @[MemPrimitives.scala 94:28:@12956.4]
  assign Mem1D_7_io_w_data_0 = _T_399[41:10]; // @[MemPrimitives.scala 95:29:@12957.4]
  assign Mem1D_7_io_w_en_0 = _T_399[42]; // @[MemPrimitives.scala 96:27:@12958.4]
  assign Mem1D_8_clock = clock; // @[:@12800.4]
  assign Mem1D_8_reset = reset; // @[:@12801.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1271[9:0]; // @[MemPrimitives.scala 131:28:@13805.4]
  assign Mem1D_8_io_r_backpressure = _T_1271[10]; // @[MemPrimitives.scala 132:32:@13806.4]
  assign Mem1D_8_io_w_ofs_0 = _T_410[9:0]; // @[MemPrimitives.scala 94:28:@12968.4]
  assign Mem1D_8_io_w_data_0 = _T_410[41:10]; // @[MemPrimitives.scala 95:29:@12969.4]
  assign Mem1D_8_io_w_en_0 = _T_410[42]; // @[MemPrimitives.scala 96:27:@12970.4]
  assign Mem1D_9_clock = clock; // @[:@12816.4]
  assign Mem1D_9_reset = reset; // @[:@12817.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1363[9:0]; // @[MemPrimitives.scala 131:28:@13894.4]
  assign Mem1D_9_io_r_backpressure = _T_1363[10]; // @[MemPrimitives.scala 132:32:@13895.4]
  assign Mem1D_9_io_w_ofs_0 = _T_421[9:0]; // @[MemPrimitives.scala 94:28:@12980.4]
  assign Mem1D_9_io_w_data_0 = _T_421[41:10]; // @[MemPrimitives.scala 95:29:@12981.4]
  assign Mem1D_9_io_w_en_0 = _T_421[42]; // @[MemPrimitives.scala 96:27:@12982.4]
  assign Mem1D_10_clock = clock; // @[:@12832.4]
  assign Mem1D_10_reset = reset; // @[:@12833.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1455[9:0]; // @[MemPrimitives.scala 131:28:@13983.4]
  assign Mem1D_10_io_r_backpressure = _T_1455[10]; // @[MemPrimitives.scala 132:32:@13984.4]
  assign Mem1D_10_io_w_ofs_0 = _T_432[9:0]; // @[MemPrimitives.scala 94:28:@12992.4]
  assign Mem1D_10_io_w_data_0 = _T_432[41:10]; // @[MemPrimitives.scala 95:29:@12993.4]
  assign Mem1D_10_io_w_en_0 = _T_432[42]; // @[MemPrimitives.scala 96:27:@12994.4]
  assign Mem1D_11_clock = clock; // @[:@12848.4]
  assign Mem1D_11_reset = reset; // @[:@12849.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1547[9:0]; // @[MemPrimitives.scala 131:28:@14072.4]
  assign Mem1D_11_io_r_backpressure = _T_1547[10]; // @[MemPrimitives.scala 132:32:@14073.4]
  assign Mem1D_11_io_w_ofs_0 = _T_443[9:0]; // @[MemPrimitives.scala 94:28:@13004.4]
  assign Mem1D_11_io_w_data_0 = _T_443[41:10]; // @[MemPrimitives.scala 95:29:@13005.4]
  assign Mem1D_11_io_w_en_0 = _T_443[42]; // @[MemPrimitives.scala 96:27:@13006.4]
  assign StickySelects_clock = clock; // @[:@13044.4]
  assign StickySelects_reset = reset; // @[:@13045.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_451; // @[MemPrimitives.scala 125:64:@13046.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_457; // @[MemPrimitives.scala 125:64:@13047.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_463; // @[MemPrimitives.scala 125:64:@13048.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_469; // @[MemPrimitives.scala 125:64:@13049.4]
  assign StickySelects_io_ins_4 = io_rPort_4_en_0 & _T_475; // @[MemPrimitives.scala 125:64:@13050.4]
  assign StickySelects_io_ins_5 = io_rPort_5_en_0 & _T_481; // @[MemPrimitives.scala 125:64:@13051.4]
  assign StickySelects_io_ins_6 = io_rPort_6_en_0 & _T_487; // @[MemPrimitives.scala 125:64:@13052.4]
  assign StickySelects_io_ins_7 = io_rPort_7_en_0 & _T_493; // @[MemPrimitives.scala 125:64:@13053.4]
  assign StickySelects_io_ins_8 = io_rPort_8_en_0 & _T_499; // @[MemPrimitives.scala 125:64:@13054.4]
  assign StickySelects_1_clock = clock; // @[:@13133.4]
  assign StickySelects_1_reset = reset; // @[:@13134.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_543; // @[MemPrimitives.scala 125:64:@13135.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_549; // @[MemPrimitives.scala 125:64:@13136.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_555; // @[MemPrimitives.scala 125:64:@13137.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_561; // @[MemPrimitives.scala 125:64:@13138.4]
  assign StickySelects_1_io_ins_4 = io_rPort_4_en_0 & _T_567; // @[MemPrimitives.scala 125:64:@13139.4]
  assign StickySelects_1_io_ins_5 = io_rPort_5_en_0 & _T_573; // @[MemPrimitives.scala 125:64:@13140.4]
  assign StickySelects_1_io_ins_6 = io_rPort_6_en_0 & _T_579; // @[MemPrimitives.scala 125:64:@13141.4]
  assign StickySelects_1_io_ins_7 = io_rPort_7_en_0 & _T_585; // @[MemPrimitives.scala 125:64:@13142.4]
  assign StickySelects_1_io_ins_8 = io_rPort_8_en_0 & _T_591; // @[MemPrimitives.scala 125:64:@13143.4]
  assign StickySelects_2_clock = clock; // @[:@13222.4]
  assign StickySelects_2_reset = reset; // @[:@13223.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@13224.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@13225.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@13226.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@13227.4]
  assign StickySelects_2_io_ins_4 = io_rPort_4_en_0 & _T_659; // @[MemPrimitives.scala 125:64:@13228.4]
  assign StickySelects_2_io_ins_5 = io_rPort_5_en_0 & _T_665; // @[MemPrimitives.scala 125:64:@13229.4]
  assign StickySelects_2_io_ins_6 = io_rPort_6_en_0 & _T_671; // @[MemPrimitives.scala 125:64:@13230.4]
  assign StickySelects_2_io_ins_7 = io_rPort_7_en_0 & _T_677; // @[MemPrimitives.scala 125:64:@13231.4]
  assign StickySelects_2_io_ins_8 = io_rPort_8_en_0 & _T_683; // @[MemPrimitives.scala 125:64:@13232.4]
  assign StickySelects_3_clock = clock; // @[:@13311.4]
  assign StickySelects_3_reset = reset; // @[:@13312.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@13313.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@13314.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@13315.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_745; // @[MemPrimitives.scala 125:64:@13316.4]
  assign StickySelects_3_io_ins_4 = io_rPort_4_en_0 & _T_751; // @[MemPrimitives.scala 125:64:@13317.4]
  assign StickySelects_3_io_ins_5 = io_rPort_5_en_0 & _T_757; // @[MemPrimitives.scala 125:64:@13318.4]
  assign StickySelects_3_io_ins_6 = io_rPort_6_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@13319.4]
  assign StickySelects_3_io_ins_7 = io_rPort_7_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@13320.4]
  assign StickySelects_3_io_ins_8 = io_rPort_8_en_0 & _T_775; // @[MemPrimitives.scala 125:64:@13321.4]
  assign StickySelects_4_clock = clock; // @[:@13400.4]
  assign StickySelects_4_reset = reset; // @[:@13401.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_819; // @[MemPrimitives.scala 125:64:@13402.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_825; // @[MemPrimitives.scala 125:64:@13403.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_831; // @[MemPrimitives.scala 125:64:@13404.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_837; // @[MemPrimitives.scala 125:64:@13405.4]
  assign StickySelects_4_io_ins_4 = io_rPort_4_en_0 & _T_843; // @[MemPrimitives.scala 125:64:@13406.4]
  assign StickySelects_4_io_ins_5 = io_rPort_5_en_0 & _T_849; // @[MemPrimitives.scala 125:64:@13407.4]
  assign StickySelects_4_io_ins_6 = io_rPort_6_en_0 & _T_855; // @[MemPrimitives.scala 125:64:@13408.4]
  assign StickySelects_4_io_ins_7 = io_rPort_7_en_0 & _T_861; // @[MemPrimitives.scala 125:64:@13409.4]
  assign StickySelects_4_io_ins_8 = io_rPort_8_en_0 & _T_867; // @[MemPrimitives.scala 125:64:@13410.4]
  assign StickySelects_5_clock = clock; // @[:@13489.4]
  assign StickySelects_5_reset = reset; // @[:@13490.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_911; // @[MemPrimitives.scala 125:64:@13491.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_917; // @[MemPrimitives.scala 125:64:@13492.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_923; // @[MemPrimitives.scala 125:64:@13493.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_929; // @[MemPrimitives.scala 125:64:@13494.4]
  assign StickySelects_5_io_ins_4 = io_rPort_4_en_0 & _T_935; // @[MemPrimitives.scala 125:64:@13495.4]
  assign StickySelects_5_io_ins_5 = io_rPort_5_en_0 & _T_941; // @[MemPrimitives.scala 125:64:@13496.4]
  assign StickySelects_5_io_ins_6 = io_rPort_6_en_0 & _T_947; // @[MemPrimitives.scala 125:64:@13497.4]
  assign StickySelects_5_io_ins_7 = io_rPort_7_en_0 & _T_953; // @[MemPrimitives.scala 125:64:@13498.4]
  assign StickySelects_5_io_ins_8 = io_rPort_8_en_0 & _T_959; // @[MemPrimitives.scala 125:64:@13499.4]
  assign StickySelects_6_clock = clock; // @[:@13578.4]
  assign StickySelects_6_reset = reset; // @[:@13579.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1003; // @[MemPrimitives.scala 125:64:@13580.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1009; // @[MemPrimitives.scala 125:64:@13581.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_1015; // @[MemPrimitives.scala 125:64:@13582.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_1021; // @[MemPrimitives.scala 125:64:@13583.4]
  assign StickySelects_6_io_ins_4 = io_rPort_4_en_0 & _T_1027; // @[MemPrimitives.scala 125:64:@13584.4]
  assign StickySelects_6_io_ins_5 = io_rPort_5_en_0 & _T_1033; // @[MemPrimitives.scala 125:64:@13585.4]
  assign StickySelects_6_io_ins_6 = io_rPort_6_en_0 & _T_1039; // @[MemPrimitives.scala 125:64:@13586.4]
  assign StickySelects_6_io_ins_7 = io_rPort_7_en_0 & _T_1045; // @[MemPrimitives.scala 125:64:@13587.4]
  assign StickySelects_6_io_ins_8 = io_rPort_8_en_0 & _T_1051; // @[MemPrimitives.scala 125:64:@13588.4]
  assign StickySelects_7_clock = clock; // @[:@13667.4]
  assign StickySelects_7_reset = reset; // @[:@13668.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1095; // @[MemPrimitives.scala 125:64:@13669.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1101; // @[MemPrimitives.scala 125:64:@13670.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1107; // @[MemPrimitives.scala 125:64:@13671.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1113; // @[MemPrimitives.scala 125:64:@13672.4]
  assign StickySelects_7_io_ins_4 = io_rPort_4_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13673.4]
  assign StickySelects_7_io_ins_5 = io_rPort_5_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13674.4]
  assign StickySelects_7_io_ins_6 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13675.4]
  assign StickySelects_7_io_ins_7 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13676.4]
  assign StickySelects_7_io_ins_8 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13677.4]
  assign StickySelects_8_clock = clock; // @[:@13756.4]
  assign StickySelects_8_reset = reset; // @[:@13757.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13758.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13759.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13760.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13761.4]
  assign StickySelects_8_io_ins_4 = io_rPort_4_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13762.4]
  assign StickySelects_8_io_ins_5 = io_rPort_5_en_0 & _T_1217; // @[MemPrimitives.scala 125:64:@13763.4]
  assign StickySelects_8_io_ins_6 = io_rPort_6_en_0 & _T_1223; // @[MemPrimitives.scala 125:64:@13764.4]
  assign StickySelects_8_io_ins_7 = io_rPort_7_en_0 & _T_1229; // @[MemPrimitives.scala 125:64:@13765.4]
  assign StickySelects_8_io_ins_8 = io_rPort_8_en_0 & _T_1235; // @[MemPrimitives.scala 125:64:@13766.4]
  assign StickySelects_9_clock = clock; // @[:@13845.4]
  assign StickySelects_9_reset = reset; // @[:@13846.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1279; // @[MemPrimitives.scala 125:64:@13847.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1285; // @[MemPrimitives.scala 125:64:@13848.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1291; // @[MemPrimitives.scala 125:64:@13849.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1297; // @[MemPrimitives.scala 125:64:@13850.4]
  assign StickySelects_9_io_ins_4 = io_rPort_4_en_0 & _T_1303; // @[MemPrimitives.scala 125:64:@13851.4]
  assign StickySelects_9_io_ins_5 = io_rPort_5_en_0 & _T_1309; // @[MemPrimitives.scala 125:64:@13852.4]
  assign StickySelects_9_io_ins_6 = io_rPort_6_en_0 & _T_1315; // @[MemPrimitives.scala 125:64:@13853.4]
  assign StickySelects_9_io_ins_7 = io_rPort_7_en_0 & _T_1321; // @[MemPrimitives.scala 125:64:@13854.4]
  assign StickySelects_9_io_ins_8 = io_rPort_8_en_0 & _T_1327; // @[MemPrimitives.scala 125:64:@13855.4]
  assign StickySelects_10_clock = clock; // @[:@13934.4]
  assign StickySelects_10_reset = reset; // @[:@13935.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1371; // @[MemPrimitives.scala 125:64:@13936.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_1377; // @[MemPrimitives.scala 125:64:@13937.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_1383; // @[MemPrimitives.scala 125:64:@13938.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_1389; // @[MemPrimitives.scala 125:64:@13939.4]
  assign StickySelects_10_io_ins_4 = io_rPort_4_en_0 & _T_1395; // @[MemPrimitives.scala 125:64:@13940.4]
  assign StickySelects_10_io_ins_5 = io_rPort_5_en_0 & _T_1401; // @[MemPrimitives.scala 125:64:@13941.4]
  assign StickySelects_10_io_ins_6 = io_rPort_6_en_0 & _T_1407; // @[MemPrimitives.scala 125:64:@13942.4]
  assign StickySelects_10_io_ins_7 = io_rPort_7_en_0 & _T_1413; // @[MemPrimitives.scala 125:64:@13943.4]
  assign StickySelects_10_io_ins_8 = io_rPort_8_en_0 & _T_1419; // @[MemPrimitives.scala 125:64:@13944.4]
  assign StickySelects_11_clock = clock; // @[:@14023.4]
  assign StickySelects_11_reset = reset; // @[:@14024.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1463; // @[MemPrimitives.scala 125:64:@14025.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1469; // @[MemPrimitives.scala 125:64:@14026.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1475; // @[MemPrimitives.scala 125:64:@14027.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1481; // @[MemPrimitives.scala 125:64:@14028.4]
  assign StickySelects_11_io_ins_4 = io_rPort_4_en_0 & _T_1487; // @[MemPrimitives.scala 125:64:@14029.4]
  assign StickySelects_11_io_ins_5 = io_rPort_5_en_0 & _T_1493; // @[MemPrimitives.scala 125:64:@14030.4]
  assign StickySelects_11_io_ins_6 = io_rPort_6_en_0 & _T_1499; // @[MemPrimitives.scala 125:64:@14031.4]
  assign StickySelects_11_io_ins_7 = io_rPort_7_en_0 & _T_1505; // @[MemPrimitives.scala 125:64:@14032.4]
  assign StickySelects_11_io_ins_8 = io_rPort_8_en_0 & _T_1511; // @[MemPrimitives.scala 125:64:@14033.4]
  assign RetimeWrapper_clock = clock; // @[:@14113.4]
  assign RetimeWrapper_reset = reset; // @[:@14114.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14116.4]
  assign RetimeWrapper_io_in = _T_451 & io_rPort_0_en_0; // @[package.scala 94:16:@14115.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14121.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14122.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14124.4]
  assign RetimeWrapper_1_io_in = _T_543 & io_rPort_0_en_0; // @[package.scala 94:16:@14123.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14129.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14130.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14132.4]
  assign RetimeWrapper_2_io_in = _T_635 & io_rPort_0_en_0; // @[package.scala 94:16:@14131.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14137.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14138.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14140.4]
  assign RetimeWrapper_3_io_in = _T_727 & io_rPort_0_en_0; // @[package.scala 94:16:@14139.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14145.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14146.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14148.4]
  assign RetimeWrapper_4_io_in = _T_819 & io_rPort_0_en_0; // @[package.scala 94:16:@14147.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14153.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14154.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14156.4]
  assign RetimeWrapper_5_io_in = _T_911 & io_rPort_0_en_0; // @[package.scala 94:16:@14155.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14161.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14162.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14164.4]
  assign RetimeWrapper_6_io_in = _T_1003 & io_rPort_0_en_0; // @[package.scala 94:16:@14163.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14169.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14170.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14172.4]
  assign RetimeWrapper_7_io_in = _T_1095 & io_rPort_0_en_0; // @[package.scala 94:16:@14171.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14177.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14178.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14180.4]
  assign RetimeWrapper_8_io_in = _T_1187 & io_rPort_0_en_0; // @[package.scala 94:16:@14179.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14185.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14186.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14188.4]
  assign RetimeWrapper_9_io_in = _T_1279 & io_rPort_0_en_0; // @[package.scala 94:16:@14187.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14193.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14194.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14196.4]
  assign RetimeWrapper_10_io_in = _T_1371 & io_rPort_0_en_0; // @[package.scala 94:16:@14195.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14201.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14202.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14204.4]
  assign RetimeWrapper_11_io_in = _T_1463 & io_rPort_0_en_0; // @[package.scala 94:16:@14203.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14257.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14258.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14260.4]
  assign RetimeWrapper_12_io_in = _T_457 & io_rPort_1_en_0; // @[package.scala 94:16:@14259.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14265.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14266.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14268.4]
  assign RetimeWrapper_13_io_in = _T_549 & io_rPort_1_en_0; // @[package.scala 94:16:@14267.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14273.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14274.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14276.4]
  assign RetimeWrapper_14_io_in = _T_641 & io_rPort_1_en_0; // @[package.scala 94:16:@14275.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14281.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14282.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14284.4]
  assign RetimeWrapper_15_io_in = _T_733 & io_rPort_1_en_0; // @[package.scala 94:16:@14283.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14289.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14290.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14292.4]
  assign RetimeWrapper_16_io_in = _T_825 & io_rPort_1_en_0; // @[package.scala 94:16:@14291.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14297.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14298.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14300.4]
  assign RetimeWrapper_17_io_in = _T_917 & io_rPort_1_en_0; // @[package.scala 94:16:@14299.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14305.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14306.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14308.4]
  assign RetimeWrapper_18_io_in = _T_1009 & io_rPort_1_en_0; // @[package.scala 94:16:@14307.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14313.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14314.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14316.4]
  assign RetimeWrapper_19_io_in = _T_1101 & io_rPort_1_en_0; // @[package.scala 94:16:@14315.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14321.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14322.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14324.4]
  assign RetimeWrapper_20_io_in = _T_1193 & io_rPort_1_en_0; // @[package.scala 94:16:@14323.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14329.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14330.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14332.4]
  assign RetimeWrapper_21_io_in = _T_1285 & io_rPort_1_en_0; // @[package.scala 94:16:@14331.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14337.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14338.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14340.4]
  assign RetimeWrapper_22_io_in = _T_1377 & io_rPort_1_en_0; // @[package.scala 94:16:@14339.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14345.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14346.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14348.4]
  assign RetimeWrapper_23_io_in = _T_1469 & io_rPort_1_en_0; // @[package.scala 94:16:@14347.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14401.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14402.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14404.4]
  assign RetimeWrapper_24_io_in = _T_463 & io_rPort_2_en_0; // @[package.scala 94:16:@14403.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14409.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14410.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14412.4]
  assign RetimeWrapper_25_io_in = _T_555 & io_rPort_2_en_0; // @[package.scala 94:16:@14411.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14417.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14418.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14420.4]
  assign RetimeWrapper_26_io_in = _T_647 & io_rPort_2_en_0; // @[package.scala 94:16:@14419.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14425.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14426.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14428.4]
  assign RetimeWrapper_27_io_in = _T_739 & io_rPort_2_en_0; // @[package.scala 94:16:@14427.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14433.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14434.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14436.4]
  assign RetimeWrapper_28_io_in = _T_831 & io_rPort_2_en_0; // @[package.scala 94:16:@14435.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14441.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14442.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14444.4]
  assign RetimeWrapper_29_io_in = _T_923 & io_rPort_2_en_0; // @[package.scala 94:16:@14443.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14449.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14450.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14452.4]
  assign RetimeWrapper_30_io_in = _T_1015 & io_rPort_2_en_0; // @[package.scala 94:16:@14451.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14457.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14458.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14460.4]
  assign RetimeWrapper_31_io_in = _T_1107 & io_rPort_2_en_0; // @[package.scala 94:16:@14459.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14465.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14466.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14468.4]
  assign RetimeWrapper_32_io_in = _T_1199 & io_rPort_2_en_0; // @[package.scala 94:16:@14467.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14473.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14474.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14476.4]
  assign RetimeWrapper_33_io_in = _T_1291 & io_rPort_2_en_0; // @[package.scala 94:16:@14475.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14481.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14482.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14484.4]
  assign RetimeWrapper_34_io_in = _T_1383 & io_rPort_2_en_0; // @[package.scala 94:16:@14483.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14489.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14490.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14492.4]
  assign RetimeWrapper_35_io_in = _T_1475 & io_rPort_2_en_0; // @[package.scala 94:16:@14491.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14545.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14546.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14548.4]
  assign RetimeWrapper_36_io_in = _T_469 & io_rPort_3_en_0; // @[package.scala 94:16:@14547.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14553.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14554.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14556.4]
  assign RetimeWrapper_37_io_in = _T_561 & io_rPort_3_en_0; // @[package.scala 94:16:@14555.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14561.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14562.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14564.4]
  assign RetimeWrapper_38_io_in = _T_653 & io_rPort_3_en_0; // @[package.scala 94:16:@14563.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14569.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14570.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14572.4]
  assign RetimeWrapper_39_io_in = _T_745 & io_rPort_3_en_0; // @[package.scala 94:16:@14571.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14577.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14578.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14580.4]
  assign RetimeWrapper_40_io_in = _T_837 & io_rPort_3_en_0; // @[package.scala 94:16:@14579.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14585.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14586.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14588.4]
  assign RetimeWrapper_41_io_in = _T_929 & io_rPort_3_en_0; // @[package.scala 94:16:@14587.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14593.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14594.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14596.4]
  assign RetimeWrapper_42_io_in = _T_1021 & io_rPort_3_en_0; // @[package.scala 94:16:@14595.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14601.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14602.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14604.4]
  assign RetimeWrapper_43_io_in = _T_1113 & io_rPort_3_en_0; // @[package.scala 94:16:@14603.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14609.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14610.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14612.4]
  assign RetimeWrapper_44_io_in = _T_1205 & io_rPort_3_en_0; // @[package.scala 94:16:@14611.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14617.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14618.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14620.4]
  assign RetimeWrapper_45_io_in = _T_1297 & io_rPort_3_en_0; // @[package.scala 94:16:@14619.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14625.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14626.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14628.4]
  assign RetimeWrapper_46_io_in = _T_1389 & io_rPort_3_en_0; // @[package.scala 94:16:@14627.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14633.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14634.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14636.4]
  assign RetimeWrapper_47_io_in = _T_1481 & io_rPort_3_en_0; // @[package.scala 94:16:@14635.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14689.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14690.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14692.4]
  assign RetimeWrapper_48_io_in = _T_475 & io_rPort_4_en_0; // @[package.scala 94:16:@14691.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14697.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14698.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14700.4]
  assign RetimeWrapper_49_io_in = _T_567 & io_rPort_4_en_0; // @[package.scala 94:16:@14699.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14705.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14706.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14708.4]
  assign RetimeWrapper_50_io_in = _T_659 & io_rPort_4_en_0; // @[package.scala 94:16:@14707.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14713.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14714.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14716.4]
  assign RetimeWrapper_51_io_in = _T_751 & io_rPort_4_en_0; // @[package.scala 94:16:@14715.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14721.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14722.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14724.4]
  assign RetimeWrapper_52_io_in = _T_843 & io_rPort_4_en_0; // @[package.scala 94:16:@14723.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14729.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14730.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14732.4]
  assign RetimeWrapper_53_io_in = _T_935 & io_rPort_4_en_0; // @[package.scala 94:16:@14731.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14737.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14738.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14740.4]
  assign RetimeWrapper_54_io_in = _T_1027 & io_rPort_4_en_0; // @[package.scala 94:16:@14739.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14745.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14746.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14748.4]
  assign RetimeWrapper_55_io_in = _T_1119 & io_rPort_4_en_0; // @[package.scala 94:16:@14747.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14753.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14754.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14756.4]
  assign RetimeWrapper_56_io_in = _T_1211 & io_rPort_4_en_0; // @[package.scala 94:16:@14755.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14761.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14762.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14764.4]
  assign RetimeWrapper_57_io_in = _T_1303 & io_rPort_4_en_0; // @[package.scala 94:16:@14763.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14769.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14770.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14772.4]
  assign RetimeWrapper_58_io_in = _T_1395 & io_rPort_4_en_0; // @[package.scala 94:16:@14771.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14777.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14778.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14780.4]
  assign RetimeWrapper_59_io_in = _T_1487 & io_rPort_4_en_0; // @[package.scala 94:16:@14779.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14833.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14834.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14836.4]
  assign RetimeWrapper_60_io_in = _T_481 & io_rPort_5_en_0; // @[package.scala 94:16:@14835.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14841.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14842.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14844.4]
  assign RetimeWrapper_61_io_in = _T_573 & io_rPort_5_en_0; // @[package.scala 94:16:@14843.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14849.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14850.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14852.4]
  assign RetimeWrapper_62_io_in = _T_665 & io_rPort_5_en_0; // @[package.scala 94:16:@14851.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14857.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14858.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14860.4]
  assign RetimeWrapper_63_io_in = _T_757 & io_rPort_5_en_0; // @[package.scala 94:16:@14859.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14865.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14866.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14868.4]
  assign RetimeWrapper_64_io_in = _T_849 & io_rPort_5_en_0; // @[package.scala 94:16:@14867.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14873.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14874.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14876.4]
  assign RetimeWrapper_65_io_in = _T_941 & io_rPort_5_en_0; // @[package.scala 94:16:@14875.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14881.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14882.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14884.4]
  assign RetimeWrapper_66_io_in = _T_1033 & io_rPort_5_en_0; // @[package.scala 94:16:@14883.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14889.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14890.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14892.4]
  assign RetimeWrapper_67_io_in = _T_1125 & io_rPort_5_en_0; // @[package.scala 94:16:@14891.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14897.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14898.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14900.4]
  assign RetimeWrapper_68_io_in = _T_1217 & io_rPort_5_en_0; // @[package.scala 94:16:@14899.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14905.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14906.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14908.4]
  assign RetimeWrapper_69_io_in = _T_1309 & io_rPort_5_en_0; // @[package.scala 94:16:@14907.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14913.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14914.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14916.4]
  assign RetimeWrapper_70_io_in = _T_1401 & io_rPort_5_en_0; // @[package.scala 94:16:@14915.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14921.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14922.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14924.4]
  assign RetimeWrapper_71_io_in = _T_1493 & io_rPort_5_en_0; // @[package.scala 94:16:@14923.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14977.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14978.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14980.4]
  assign RetimeWrapper_72_io_in = _T_487 & io_rPort_6_en_0; // @[package.scala 94:16:@14979.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14985.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14986.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14988.4]
  assign RetimeWrapper_73_io_in = _T_579 & io_rPort_6_en_0; // @[package.scala 94:16:@14987.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14993.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14994.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14996.4]
  assign RetimeWrapper_74_io_in = _T_671 & io_rPort_6_en_0; // @[package.scala 94:16:@14995.4]
  assign RetimeWrapper_75_clock = clock; // @[:@15001.4]
  assign RetimeWrapper_75_reset = reset; // @[:@15002.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15004.4]
  assign RetimeWrapper_75_io_in = _T_763 & io_rPort_6_en_0; // @[package.scala 94:16:@15003.4]
  assign RetimeWrapper_76_clock = clock; // @[:@15009.4]
  assign RetimeWrapper_76_reset = reset; // @[:@15010.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15012.4]
  assign RetimeWrapper_76_io_in = _T_855 & io_rPort_6_en_0; // @[package.scala 94:16:@15011.4]
  assign RetimeWrapper_77_clock = clock; // @[:@15017.4]
  assign RetimeWrapper_77_reset = reset; // @[:@15018.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15020.4]
  assign RetimeWrapper_77_io_in = _T_947 & io_rPort_6_en_0; // @[package.scala 94:16:@15019.4]
  assign RetimeWrapper_78_clock = clock; // @[:@15025.4]
  assign RetimeWrapper_78_reset = reset; // @[:@15026.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15028.4]
  assign RetimeWrapper_78_io_in = _T_1039 & io_rPort_6_en_0; // @[package.scala 94:16:@15027.4]
  assign RetimeWrapper_79_clock = clock; // @[:@15033.4]
  assign RetimeWrapper_79_reset = reset; // @[:@15034.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15036.4]
  assign RetimeWrapper_79_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@15035.4]
  assign RetimeWrapper_80_clock = clock; // @[:@15041.4]
  assign RetimeWrapper_80_reset = reset; // @[:@15042.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15044.4]
  assign RetimeWrapper_80_io_in = _T_1223 & io_rPort_6_en_0; // @[package.scala 94:16:@15043.4]
  assign RetimeWrapper_81_clock = clock; // @[:@15049.4]
  assign RetimeWrapper_81_reset = reset; // @[:@15050.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15052.4]
  assign RetimeWrapper_81_io_in = _T_1315 & io_rPort_6_en_0; // @[package.scala 94:16:@15051.4]
  assign RetimeWrapper_82_clock = clock; // @[:@15057.4]
  assign RetimeWrapper_82_reset = reset; // @[:@15058.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15060.4]
  assign RetimeWrapper_82_io_in = _T_1407 & io_rPort_6_en_0; // @[package.scala 94:16:@15059.4]
  assign RetimeWrapper_83_clock = clock; // @[:@15065.4]
  assign RetimeWrapper_83_reset = reset; // @[:@15066.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15068.4]
  assign RetimeWrapper_83_io_in = _T_1499 & io_rPort_6_en_0; // @[package.scala 94:16:@15067.4]
  assign RetimeWrapper_84_clock = clock; // @[:@15121.4]
  assign RetimeWrapper_84_reset = reset; // @[:@15122.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15124.4]
  assign RetimeWrapper_84_io_in = _T_493 & io_rPort_7_en_0; // @[package.scala 94:16:@15123.4]
  assign RetimeWrapper_85_clock = clock; // @[:@15129.4]
  assign RetimeWrapper_85_reset = reset; // @[:@15130.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15132.4]
  assign RetimeWrapper_85_io_in = _T_585 & io_rPort_7_en_0; // @[package.scala 94:16:@15131.4]
  assign RetimeWrapper_86_clock = clock; // @[:@15137.4]
  assign RetimeWrapper_86_reset = reset; // @[:@15138.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15140.4]
  assign RetimeWrapper_86_io_in = _T_677 & io_rPort_7_en_0; // @[package.scala 94:16:@15139.4]
  assign RetimeWrapper_87_clock = clock; // @[:@15145.4]
  assign RetimeWrapper_87_reset = reset; // @[:@15146.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15148.4]
  assign RetimeWrapper_87_io_in = _T_769 & io_rPort_7_en_0; // @[package.scala 94:16:@15147.4]
  assign RetimeWrapper_88_clock = clock; // @[:@15153.4]
  assign RetimeWrapper_88_reset = reset; // @[:@15154.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15156.4]
  assign RetimeWrapper_88_io_in = _T_861 & io_rPort_7_en_0; // @[package.scala 94:16:@15155.4]
  assign RetimeWrapper_89_clock = clock; // @[:@15161.4]
  assign RetimeWrapper_89_reset = reset; // @[:@15162.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15164.4]
  assign RetimeWrapper_89_io_in = _T_953 & io_rPort_7_en_0; // @[package.scala 94:16:@15163.4]
  assign RetimeWrapper_90_clock = clock; // @[:@15169.4]
  assign RetimeWrapper_90_reset = reset; // @[:@15170.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15172.4]
  assign RetimeWrapper_90_io_in = _T_1045 & io_rPort_7_en_0; // @[package.scala 94:16:@15171.4]
  assign RetimeWrapper_91_clock = clock; // @[:@15177.4]
  assign RetimeWrapper_91_reset = reset; // @[:@15178.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15180.4]
  assign RetimeWrapper_91_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@15179.4]
  assign RetimeWrapper_92_clock = clock; // @[:@15185.4]
  assign RetimeWrapper_92_reset = reset; // @[:@15186.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15188.4]
  assign RetimeWrapper_92_io_in = _T_1229 & io_rPort_7_en_0; // @[package.scala 94:16:@15187.4]
  assign RetimeWrapper_93_clock = clock; // @[:@15193.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15194.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15196.4]
  assign RetimeWrapper_93_io_in = _T_1321 & io_rPort_7_en_0; // @[package.scala 94:16:@15195.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15201.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15202.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15204.4]
  assign RetimeWrapper_94_io_in = _T_1413 & io_rPort_7_en_0; // @[package.scala 94:16:@15203.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15209.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15210.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15212.4]
  assign RetimeWrapper_95_io_in = _T_1505 & io_rPort_7_en_0; // @[package.scala 94:16:@15211.4]
  assign RetimeWrapper_96_clock = clock; // @[:@15265.4]
  assign RetimeWrapper_96_reset = reset; // @[:@15266.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15268.4]
  assign RetimeWrapper_96_io_in = _T_499 & io_rPort_8_en_0; // @[package.scala 94:16:@15267.4]
  assign RetimeWrapper_97_clock = clock; // @[:@15273.4]
  assign RetimeWrapper_97_reset = reset; // @[:@15274.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15276.4]
  assign RetimeWrapper_97_io_in = _T_591 & io_rPort_8_en_0; // @[package.scala 94:16:@15275.4]
  assign RetimeWrapper_98_clock = clock; // @[:@15281.4]
  assign RetimeWrapper_98_reset = reset; // @[:@15282.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15284.4]
  assign RetimeWrapper_98_io_in = _T_683 & io_rPort_8_en_0; // @[package.scala 94:16:@15283.4]
  assign RetimeWrapper_99_clock = clock; // @[:@15289.4]
  assign RetimeWrapper_99_reset = reset; // @[:@15290.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15292.4]
  assign RetimeWrapper_99_io_in = _T_775 & io_rPort_8_en_0; // @[package.scala 94:16:@15291.4]
  assign RetimeWrapper_100_clock = clock; // @[:@15297.4]
  assign RetimeWrapper_100_reset = reset; // @[:@15298.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15300.4]
  assign RetimeWrapper_100_io_in = _T_867 & io_rPort_8_en_0; // @[package.scala 94:16:@15299.4]
  assign RetimeWrapper_101_clock = clock; // @[:@15305.4]
  assign RetimeWrapper_101_reset = reset; // @[:@15306.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15308.4]
  assign RetimeWrapper_101_io_in = _T_959 & io_rPort_8_en_0; // @[package.scala 94:16:@15307.4]
  assign RetimeWrapper_102_clock = clock; // @[:@15313.4]
  assign RetimeWrapper_102_reset = reset; // @[:@15314.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15316.4]
  assign RetimeWrapper_102_io_in = _T_1051 & io_rPort_8_en_0; // @[package.scala 94:16:@15315.4]
  assign RetimeWrapper_103_clock = clock; // @[:@15321.4]
  assign RetimeWrapper_103_reset = reset; // @[:@15322.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15324.4]
  assign RetimeWrapper_103_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@15323.4]
  assign RetimeWrapper_104_clock = clock; // @[:@15329.4]
  assign RetimeWrapper_104_reset = reset; // @[:@15330.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15332.4]
  assign RetimeWrapper_104_io_in = _T_1235 & io_rPort_8_en_0; // @[package.scala 94:16:@15331.4]
  assign RetimeWrapper_105_clock = clock; // @[:@15337.4]
  assign RetimeWrapper_105_reset = reset; // @[:@15338.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15340.4]
  assign RetimeWrapper_105_io_in = _T_1327 & io_rPort_8_en_0; // @[package.scala 94:16:@15339.4]
  assign RetimeWrapper_106_clock = clock; // @[:@15345.4]
  assign RetimeWrapper_106_reset = reset; // @[:@15346.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15348.4]
  assign RetimeWrapper_106_io_in = _T_1419 & io_rPort_8_en_0; // @[package.scala 94:16:@15347.4]
  assign RetimeWrapper_107_clock = clock; // @[:@15353.4]
  assign RetimeWrapper_107_reset = reset; // @[:@15354.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15356.4]
  assign RetimeWrapper_107_io_in = _T_1511 & io_rPort_8_en_0; // @[package.scala 94:16:@15355.4]
endmodule
module Divider( // @[:@16978.2]
  input         clock, // @[:@16979.4]
  input         io_flow, // @[:@16981.4]
  input  [31:0] io_dividend, // @[:@16981.4]
  input  [31:0] io_divisor, // @[:@16981.4]
  output [31:0] io_out // @[:@16981.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire [29:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@16999.4]
  div_32_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@16983.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[31:2]; // @[ZynqBlackBoxes.scala 34:37:@16999.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@17000.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@16997.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@16996.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@16995.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@16994.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@16993.4 ZynqBlackBoxes.scala 33:17:@16998.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@16992.4]
endmodule
module x235_div( // @[:@17038.2]
  input         clock, // @[:@17039.4]
  input  [31:0] io_a, // @[:@17041.4]
  input         io_flow, // @[:@17041.4]
  output [31:0] io_result // @[:@17041.4]
);
  wire  x235_div_clock; // @[BigIPZynq.scala 25:21:@17049.4]
  wire  x235_div_io_flow; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] x235_div_io_dividend; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] x235_div_io_divisor; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] x235_div_io_out; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@17062.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@17062.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@17047.4]
  wire [31:0] _T_19; // @[BigIPZynq.scala 29:16:@17057.4]
  Divider x235_div ( // @[BigIPZynq.scala 25:21:@17049.4]
    .clock(x235_div_clock),
    .io_flow(x235_div_io_flow),
    .io_dividend(x235_div_io_dividend),
    .io_divisor(x235_div_io_divisor),
    .io_out(x235_div_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@17062.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@17047.4]
  assign _T_19 = $signed(x235_div_io_out); // @[BigIPZynq.scala 29:16:@17057.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@17070.4]
  assign x235_div_clock = clock; // @[:@17050.4]
  assign x235_div_io_flow = io_flow; // @[BigIPZynq.scala 28:17:@17056.4]
  assign x235_div_io_dividend = $unsigned(_T_15); // @[BigIPZynq.scala 26:21:@17053.4]
  assign x235_div_io_divisor = 32'h3; // @[BigIPZynq.scala 27:20:@17055.4]
  assign __io_b = $unsigned(_T_19); // @[Math.scala 721:17:@17065.4]
endmodule
module RetimeWrapper_184( // @[:@17084.2]
  input         clock, // @[:@17085.4]
  input         reset, // @[:@17086.4]
  input         io_flow, // @[:@17087.4]
  input  [31:0] io_in, // @[:@17087.4]
  output [31:0] io_out // @[:@17087.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@17089.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17102.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17101.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17100.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17099.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17098.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17096.4]
endmodule
module RetimeWrapper_186( // @[:@17295.2]
  input         clock, // @[:@17296.4]
  input         reset, // @[:@17297.4]
  input         io_flow, // @[:@17298.4]
  input  [31:0] io_in, // @[:@17298.4]
  output [31:0] io_out // @[:@17298.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@17300.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17313.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17312.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17311.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17310.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17309.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17307.4]
endmodule
module RetimeWrapper_187( // @[:@17327.2]
  input   clock, // @[:@17328.4]
  input   reset, // @[:@17329.4]
  input   io_flow, // @[:@17330.4]
  input   io_in, // @[:@17330.4]
  output  io_out // @[:@17330.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@17332.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17345.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17344.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@17343.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17342.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17341.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17339.4]
endmodule
module RetimeWrapper_188( // @[:@17359.2]
  input         clock, // @[:@17360.4]
  input         reset, // @[:@17361.4]
  input         io_flow, // @[:@17362.4]
  input  [31:0] io_in, // @[:@17362.4]
  output [31:0] io_out // @[:@17362.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@17364.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17377.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17376.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17375.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17374.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17373.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17371.4]
endmodule
module RetimeWrapper_190( // @[:@17423.2]
  input         clock, // @[:@17424.4]
  input         reset, // @[:@17425.4]
  input         io_flow, // @[:@17426.4]
  input  [31:0] io_in, // @[:@17426.4]
  output [31:0] io_out // @[:@17426.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17428.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17428.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17428.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17428.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17428.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17428.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@17428.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17441.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17440.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17439.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17438.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17437.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17435.4]
endmodule
module RetimeWrapper_192( // @[:@17487.2]
  input         clock, // @[:@17488.4]
  input         reset, // @[:@17489.4]
  input         io_flow, // @[:@17490.4]
  input  [31:0] io_in, // @[:@17490.4]
  output [31:0] io_out // @[:@17490.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@17492.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17505.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17504.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17503.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17502.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17501.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17499.4]
endmodule
module RetimeWrapper_196( // @[:@17615.2]
  input         clock, // @[:@17616.4]
  input         reset, // @[:@17617.4]
  input         io_flow, // @[:@17618.4]
  input  [31:0] io_in, // @[:@17618.4]
  output [31:0] io_out // @[:@17618.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(37)) sr ( // @[RetimeShiftRegister.scala 15:20:@17620.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17633.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17632.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17631.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17630.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17629.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17627.4]
endmodule
module RetimeWrapper_197( // @[:@17647.2]
  input   clock, // @[:@17648.4]
  input   reset, // @[:@17649.4]
  input   io_flow, // @[:@17650.4]
  input   io_in, // @[:@17650.4]
  output  io_out // @[:@17650.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@17652.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17665.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17664.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@17663.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17662.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17661.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17659.4]
endmodule
module RetimeWrapper_198( // @[:@17679.2]
  input         clock, // @[:@17680.4]
  input         reset, // @[:@17681.4]
  input         io_flow, // @[:@17682.4]
  input  [31:0] io_in, // @[:@17682.4]
  output [31:0] io_out // @[:@17682.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@17684.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17697.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17696.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17695.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17694.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17693.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17691.4]
endmodule
module RetimeWrapper_201( // @[:@17775.2]
  input         clock, // @[:@17776.4]
  input         reset, // @[:@17777.4]
  input         io_flow, // @[:@17778.4]
  input  [31:0] io_in, // @[:@17778.4]
  output [31:0] io_out // @[:@17778.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17780.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17780.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17780.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17780.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17780.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17780.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@17780.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17793.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17792.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17791.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17790.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17789.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17787.4]
endmodule
module RetimeWrapper_218( // @[:@19604.2]
  input         clock, // @[:@19605.4]
  input         reset, // @[:@19606.4]
  input         io_flow, // @[:@19607.4]
  input  [31:0] io_in, // @[:@19607.4]
  output [31:0] io_out // @[:@19607.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(43)) sr ( // @[RetimeShiftRegister.scala 15:20:@19609.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@19622.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@19621.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@19620.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@19619.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@19618.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@19616.4]
endmodule
module RetimeWrapper_220( // @[:@19815.2]
  input   clock, // @[:@19816.4]
  input   reset, // @[:@19817.4]
  input   io_flow, // @[:@19818.4]
  input   io_in, // @[:@19818.4]
  output  io_out // @[:@19818.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@19820.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@19833.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@19832.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@19831.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@19830.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@19829.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@19827.4]
endmodule
module RetimeWrapper_247( // @[:@22406.2]
  input         clock, // @[:@22407.4]
  input         reset, // @[:@22408.4]
  input         io_flow, // @[:@22409.4]
  input  [31:0] io_in, // @[:@22409.4]
  output [31:0] io_out // @[:@22409.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22411.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22411.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22411.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22411.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22411.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22411.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@22411.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22424.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22423.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22422.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22421.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22420.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22418.4]
endmodule
module RetimeWrapper_254( // @[:@22777.2]
  input         clock, // @[:@22778.4]
  input         reset, // @[:@22779.4]
  input         io_flow, // @[:@22780.4]
  input  [31:0] io_in, // @[:@22780.4]
  output [31:0] io_out // @[:@22780.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@22782.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22795.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22794.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22793.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22792.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22791.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22789.4]
endmodule
module Multiplier( // @[:@24605.2]
  input         clock, // @[:@24606.4]
  input         io_flow, // @[:@24608.4]
  input  [31:0] io_a, // @[:@24608.4]
  input  [31:0] io_b, // @[:@24608.4]
  output [31:0] io_out // @[:@24608.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@24610.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@24620.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@24618.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@24617.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@24619.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@24616.4]
endmodule
module x305( // @[:@24640.2]
  input         clock, // @[:@24641.4]
  input  [31:0] io_a, // @[:@24643.4]
  input  [31:0] io_b, // @[:@24643.4]
  input         io_flow, // @[:@24643.4]
  output [31:0] io_result // @[:@24643.4]
);
  wire  x305_clock; // @[BigIPZynq.scala 63:21:@24650.4]
  wire  x305_io_flow; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] x305_io_a; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] x305_io_b; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] x305_io_out; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@24659.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@24659.4]
  Multiplier x305 ( // @[BigIPZynq.scala 63:21:@24650.4]
    .clock(x305_clock),
    .io_flow(x305_io_flow),
    .io_a(x305_io_a),
    .io_b(x305_io_b),
    .io_out(x305_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@24659.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@24667.4]
  assign x305_clock = clock; // @[:@24651.4]
  assign x305_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@24655.4]
  assign x305_io_a = io_a; // @[BigIPZynq.scala 64:14:@24653.4]
  assign x305_io_b = io_b; // @[BigIPZynq.scala 65:14:@24654.4]
  assign fix2fixBox_io_a = x305_io_out; // @[Math.scala 254:23:@24662.4]
endmodule
module fix2fixBox_140( // @[:@25261.2]
  input  [31:0] io_a, // @[:@25264.4]
  output [32:0] io_b // @[:@25264.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@25278.4]
endmodule
module __89( // @[:@25280.2]
  input  [31:0] io_b, // @[:@25283.4]
  output [32:0] io_result // @[:@25283.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@25288.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@25288.4]
  fix2fixBox_140 fix2fixBox ( // @[BigIPZynq.scala 219:30:@25288.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@25296.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@25291.4]
endmodule
module x314_x13( // @[:@25392.2]
  input         clock, // @[:@25393.4]
  input         reset, // @[:@25394.4]
  input  [31:0] io_a, // @[:@25395.4]
  input  [31:0] io_b, // @[:@25395.4]
  input         io_flow, // @[:@25395.4]
  output [31:0] io_result // @[:@25395.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@25403.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@25403.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@25410.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@25410.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@25420.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@25420.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@25420.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@25420.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@25420.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@25408.4 Math.scala 724:14:@25409.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@25415.4 Math.scala 724:14:@25416.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@25417.4]
  __89 _ ( // @[Math.scala 720:24:@25403.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __89 __1 ( // @[Math.scala 720:24:@25410.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@25420.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@25408.4 Math.scala 724:14:@25409.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@25415.4 Math.scala 724:14:@25416.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@25417.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@25428.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@25406.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@25413.4]
  assign fix2fixBox_clock = clock; // @[:@25421.4]
  assign fix2fixBox_reset = reset; // @[:@25422.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@25423.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@25426.4]
endmodule
module RetimeWrapper_286( // @[:@26456.2]
  input         clock, // @[:@26457.4]
  input         reset, // @[:@26458.4]
  input         io_flow, // @[:@26459.4]
  input  [31:0] io_in, // @[:@26459.4]
  output [31:0] io_out // @[:@26459.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26461.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26474.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26473.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26472.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26471.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26470.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26468.4]
endmodule
module fix2fixBox_164( // @[:@26645.2]
  input  [31:0] io_a, // @[:@26648.4]
  output [31:0] io_b // @[:@26648.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@26658.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@26658.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@26661.4]
endmodule
module x322( // @[:@26663.2]
  input  [31:0] io_b, // @[:@26666.4]
  output [31:0] io_result // @[:@26666.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@26671.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@26671.4]
  fix2fixBox_164 fix2fixBox ( // @[BigIPZynq.scala 219:30:@26671.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@26679.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@26674.4]
endmodule
module Multiplier_9( // @[:@26691.2]
  input         clock, // @[:@26692.4]
  input         io_flow, // @[:@26694.4]
  input  [38:0] io_a, // @[:@26694.4]
  input  [38:0] io_b, // @[:@26694.4]
  output [38:0] io_out // @[:@26694.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@26696.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@26706.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@26704.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@26703.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@26705.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@26702.4]
endmodule
module fix2fixBox_165( // @[:@26708.2]
  input  [38:0] io_a, // @[:@26711.4]
  output [31:0] io_b // @[:@26711.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@26719.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@26722.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@26719.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@26722.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@26725.4]
endmodule
module x323_mul( // @[:@26727.2]
  input         clock, // @[:@26728.4]
  input  [31:0] io_a, // @[:@26730.4]
  input  [31:0] io_b, // @[:@26730.4]
  input         io_flow, // @[:@26730.4]
  output [31:0] io_result // @[:@26730.4]
);
  wire  x323_mul_clock; // @[BigIPZynq.scala 63:21:@26745.4]
  wire  x323_mul_io_flow; // @[BigIPZynq.scala 63:21:@26745.4]
  wire [38:0] x323_mul_io_a; // @[BigIPZynq.scala 63:21:@26745.4]
  wire [38:0] x323_mul_io_b; // @[BigIPZynq.scala 63:21:@26745.4]
  wire [38:0] x323_mul_io_out; // @[BigIPZynq.scala 63:21:@26745.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@26753.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@26753.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@26737.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@26739.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@26741.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@26743.4]
  Multiplier_9 x323_mul ( // @[BigIPZynq.scala 63:21:@26745.4]
    .clock(x323_mul_clock),
    .io_flow(x323_mul_io_flow),
    .io_a(x323_mul_io_a),
    .io_b(x323_mul_io_b),
    .io_out(x323_mul_io_out)
  );
  fix2fixBox_165 fix2fixBox ( // @[Math.scala 253:30:@26753.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@26737.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@26739.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@26741.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@26743.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@26761.4]
  assign x323_mul_clock = clock; // @[:@26746.4]
  assign x323_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@26750.4]
  assign x323_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@26748.4]
  assign x323_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@26749.4]
  assign fix2fixBox_io_a = x323_mul_io_out; // @[Math.scala 254:23:@26756.4]
endmodule
module fix2fixBox_166( // @[:@26763.2]
  input  [31:0] io_a, // @[:@26766.4]
  output [31:0] io_b // @[:@26766.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@26778.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@26778.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@26781.4]
endmodule
module x324( // @[:@26783.2]
  input  [31:0] io_b, // @[:@26786.4]
  output [31:0] io_result // @[:@26786.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@26791.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@26791.4]
  fix2fixBox_166 fix2fixBox ( // @[BigIPZynq.scala 219:30:@26791.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@26799.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@26794.4]
endmodule
module RetimeWrapper_288( // @[:@26813.2]
  input         clock, // @[:@26814.4]
  input         reset, // @[:@26815.4]
  input         io_flow, // @[:@26816.4]
  input  [31:0] io_in, // @[:@26816.4]
  output [31:0] io_out // @[:@26816.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26818.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26818.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26818.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26818.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26818.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26818.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@26818.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26831.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26830.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26829.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26828.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26827.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26825.4]
endmodule
module x325_sub( // @[:@26964.2]
  input         clock, // @[:@26965.4]
  input         reset, // @[:@26966.4]
  input  [31:0] io_a, // @[:@26967.4]
  input  [31:0] io_b, // @[:@26967.4]
  input         io_flow, // @[:@26967.4]
  output [31:0] io_result // @[:@26967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@26975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@26975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@26982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@26982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@26993.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@26993.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@26993.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@26993.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@26993.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@26980.4 Math.scala 724:14:@26981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@26987.4 Math.scala 724:14:@26988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@26989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@26990.4]
  __89 _ ( // @[Math.scala 720:24:@26975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __89 __1 ( // @[Math.scala 720:24:@26982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@26993.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@26980.4 Math.scala 724:14:@26981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@26987.4 Math.scala 724:14:@26988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@26989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@26990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@27001.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@26978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@26985.4]
  assign fix2fixBox_clock = clock; // @[:@26994.4]
  assign fix2fixBox_reset = reset; // @[:@26995.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@26996.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@26999.4]
endmodule
module x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@27754.2]
  input          clock, // @[:@27755.4]
  input          reset, // @[:@27756.4]
  output         io_in_x194_TREADY, // @[:@27757.4]
  input  [255:0] io_in_x194_TDATA, // @[:@27757.4]
  input  [7:0]   io_in_x194_TID, // @[:@27757.4]
  input  [7:0]   io_in_x194_TDEST, // @[:@27757.4]
  output         io_in_x195_TVALID, // @[:@27757.4]
  input          io_in_x195_TREADY, // @[:@27757.4]
  output [255:0] io_in_x195_TDATA, // @[:@27757.4]
  input          io_sigsIn_backpressure, // @[:@27757.4]
  input          io_sigsIn_datapathEn, // @[:@27757.4]
  input          io_sigsIn_break, // @[:@27757.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@27757.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@27757.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@27757.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@27757.4]
  input          io_rr // @[:@27757.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@27771.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@27771.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@27783.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@27783.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@27806.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@27806.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@27806.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@27806.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@27806.4]
  wire  x227_lb_0_clock; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_reset; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_8_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_8_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_8_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_8_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_8_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_8_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_7_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_7_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_7_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_7_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_7_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_7_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_6_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_6_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_6_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_6_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_6_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_6_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_5_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_5_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_5_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_5_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_5_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_5_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_4_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_4_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_4_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_4_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_4_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_4_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_3_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_3_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_3_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_3_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_3_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_3_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_2_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_2_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_2_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_2_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_2_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_2_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_1_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_1_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_1_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_1_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_1_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_1_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_rPort_0_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_rPort_0_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_rPort_0_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_0_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_rPort_0_backpressure; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_rPort_0_output_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [1:0] x227_lb_0_io_wPort_0_banks_1; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [2:0] x227_lb_0_io_wPort_0_banks_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [9:0] x227_lb_0_io_wPort_0_ofs_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire [31:0] x227_lb_0_io_wPort_0_data_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x227_lb_0_io_wPort_0_en_0; // @[m_x227_lb_0.scala 35:17:@27816.4]
  wire  x398_sum_1_clock; // @[Math.scala 150:24:@27941.4]
  wire  x398_sum_1_reset; // @[Math.scala 150:24:@27941.4]
  wire [31:0] x398_sum_1_io_a; // @[Math.scala 150:24:@27941.4]
  wire [31:0] x398_sum_1_io_b; // @[Math.scala 150:24:@27941.4]
  wire  x398_sum_1_io_flow; // @[Math.scala 150:24:@27941.4]
  wire [31:0] x398_sum_1_io_result; // @[Math.scala 150:24:@27941.4]
  wire  x401_sum_1_clock; // @[Math.scala 150:24:@27979.4]
  wire  x401_sum_1_reset; // @[Math.scala 150:24:@27979.4]
  wire [31:0] x401_sum_1_io_a; // @[Math.scala 150:24:@27979.4]
  wire [31:0] x401_sum_1_io_b; // @[Math.scala 150:24:@27979.4]
  wire  x401_sum_1_io_flow; // @[Math.scala 150:24:@27979.4]
  wire [31:0] x401_sum_1_io_result; // @[Math.scala 150:24:@27979.4]
  wire  x404_sum_1_clock; // @[Math.scala 150:24:@28017.4]
  wire  x404_sum_1_reset; // @[Math.scala 150:24:@28017.4]
  wire [31:0] x404_sum_1_io_a; // @[Math.scala 150:24:@28017.4]
  wire [31:0] x404_sum_1_io_b; // @[Math.scala 150:24:@28017.4]
  wire  x404_sum_1_io_flow; // @[Math.scala 150:24:@28017.4]
  wire [31:0] x404_sum_1_io_result; // @[Math.scala 150:24:@28017.4]
  wire  x407_sum_1_clock; // @[Math.scala 150:24:@28055.4]
  wire  x407_sum_1_reset; // @[Math.scala 150:24:@28055.4]
  wire [31:0] x407_sum_1_io_a; // @[Math.scala 150:24:@28055.4]
  wire [31:0] x407_sum_1_io_b; // @[Math.scala 150:24:@28055.4]
  wire  x407_sum_1_io_flow; // @[Math.scala 150:24:@28055.4]
  wire [31:0] x407_sum_1_io_result; // @[Math.scala 150:24:@28055.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@28078.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@28078.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@28078.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@28078.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@28078.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@28096.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@28096.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@28096.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@28096.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@28096.4]
  wire  x410_sum_1_clock; // @[Math.scala 150:24:@28109.4]
  wire  x410_sum_1_reset; // @[Math.scala 150:24:@28109.4]
  wire [31:0] x410_sum_1_io_a; // @[Math.scala 150:24:@28109.4]
  wire [31:0] x410_sum_1_io_b; // @[Math.scala 150:24:@28109.4]
  wire  x410_sum_1_io_flow; // @[Math.scala 150:24:@28109.4]
  wire [31:0] x410_sum_1_io_result; // @[Math.scala 150:24:@28109.4]
  wire  x413_sum_1_clock; // @[Math.scala 150:24:@28147.4]
  wire  x413_sum_1_reset; // @[Math.scala 150:24:@28147.4]
  wire [31:0] x413_sum_1_io_a; // @[Math.scala 150:24:@28147.4]
  wire [31:0] x413_sum_1_io_b; // @[Math.scala 150:24:@28147.4]
  wire  x413_sum_1_io_flow; // @[Math.scala 150:24:@28147.4]
  wire [31:0] x413_sum_1_io_result; // @[Math.scala 150:24:@28147.4]
  wire  x416_sub_1_clock; // @[Math.scala 191:24:@28173.4]
  wire  x416_sub_1_reset; // @[Math.scala 191:24:@28173.4]
  wire [31:0] x416_sub_1_io_a; // @[Math.scala 191:24:@28173.4]
  wire [31:0] x416_sub_1_io_b; // @[Math.scala 191:24:@28173.4]
  wire  x416_sub_1_io_flow; // @[Math.scala 191:24:@28173.4]
  wire [31:0] x416_sub_1_io_result; // @[Math.scala 191:24:@28173.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@28183.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@28183.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@28183.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@28183.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@28183.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@28192.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@28192.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@28192.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@28192.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@28192.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@28201.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@28201.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@28201.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@28201.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@28201.4]
  wire  x420_sum_1_clock; // @[Math.scala 150:24:@28240.4]
  wire  x420_sum_1_reset; // @[Math.scala 150:24:@28240.4]
  wire [31:0] x420_sum_1_io_a; // @[Math.scala 150:24:@28240.4]
  wire [31:0] x420_sum_1_io_b; // @[Math.scala 150:24:@28240.4]
  wire  x420_sum_1_io_flow; // @[Math.scala 150:24:@28240.4]
  wire [31:0] x420_sum_1_io_result; // @[Math.scala 150:24:@28240.4]
  wire  x235_div_1_clock; // @[Math.scala 327:24:@28252.4]
  wire [31:0] x235_div_1_io_a; // @[Math.scala 327:24:@28252.4]
  wire  x235_div_1_io_flow; // @[Math.scala 327:24:@28252.4]
  wire [31:0] x235_div_1_io_result; // @[Math.scala 327:24:@28252.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@28262.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@28262.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@28262.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@28262.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@28262.4]
  wire  x236_sum_1_clock; // @[Math.scala 150:24:@28271.4]
  wire  x236_sum_1_reset; // @[Math.scala 150:24:@28271.4]
  wire [31:0] x236_sum_1_io_a; // @[Math.scala 150:24:@28271.4]
  wire [31:0] x236_sum_1_io_b; // @[Math.scala 150:24:@28271.4]
  wire  x236_sum_1_io_flow; // @[Math.scala 150:24:@28271.4]
  wire [31:0] x236_sum_1_io_result; // @[Math.scala 150:24:@28271.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@28281.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@28281.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@28281.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@28281.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@28281.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@28290.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@28290.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@28290.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@28290.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@28290.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@28299.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@28299.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@28299.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@28299.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@28299.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@28308.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@28308.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@28308.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@28308.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@28308.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@28317.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@28317.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@28317.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@28317.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@28317.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@28328.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@28328.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@28328.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@28328.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@28328.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@28349.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@28349.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@28372.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@28372.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@28372.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@28372.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@28372.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@28388.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@28403.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@28403.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@28403.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@28403.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@28403.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@28412.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@28412.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@28412.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@28412.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@28412.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@28421.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@28421.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@28421.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@28421.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@28421.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@28430.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@28430.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@28430.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@28430.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@28430.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@28448.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@28448.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@28448.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@28448.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@28448.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@28460.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@28460.4]
  wire  x245_rdcol_1_clock; // @[Math.scala 191:24:@28483.4]
  wire  x245_rdcol_1_reset; // @[Math.scala 191:24:@28483.4]
  wire [31:0] x245_rdcol_1_io_a; // @[Math.scala 191:24:@28483.4]
  wire [31:0] x245_rdcol_1_io_b; // @[Math.scala 191:24:@28483.4]
  wire  x245_rdcol_1_io_flow; // @[Math.scala 191:24:@28483.4]
  wire [31:0] x245_rdcol_1_io_result; // @[Math.scala 191:24:@28483.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@28498.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@28498.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@28498.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@28498.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@28498.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@28507.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@28507.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@28507.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@28507.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@28507.4]
  wire  x423_sum_1_clock; // @[Math.scala 150:24:@28550.4]
  wire  x423_sum_1_reset; // @[Math.scala 150:24:@28550.4]
  wire [31:0] x423_sum_1_io_a; // @[Math.scala 150:24:@28550.4]
  wire [31:0] x423_sum_1_io_b; // @[Math.scala 150:24:@28550.4]
  wire  x423_sum_1_io_flow; // @[Math.scala 150:24:@28550.4]
  wire [31:0] x423_sum_1_io_result; // @[Math.scala 150:24:@28550.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@28573.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@28573.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@28573.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@28573.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@28573.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@28591.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@28591.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@28591.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@28591.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@28591.4]
  wire  x426_sum_1_clock; // @[Math.scala 150:24:@28604.4]
  wire  x426_sum_1_reset; // @[Math.scala 150:24:@28604.4]
  wire [31:0] x426_sum_1_io_a; // @[Math.scala 150:24:@28604.4]
  wire [31:0] x426_sum_1_io_b; // @[Math.scala 150:24:@28604.4]
  wire  x426_sum_1_io_flow; // @[Math.scala 150:24:@28604.4]
  wire [31:0] x426_sum_1_io_result; // @[Math.scala 150:24:@28604.4]
  wire  x429_sum_1_clock; // @[Math.scala 150:24:@28642.4]
  wire  x429_sum_1_reset; // @[Math.scala 150:24:@28642.4]
  wire [31:0] x429_sum_1_io_a; // @[Math.scala 150:24:@28642.4]
  wire [31:0] x429_sum_1_io_b; // @[Math.scala 150:24:@28642.4]
  wire  x429_sum_1_io_flow; // @[Math.scala 150:24:@28642.4]
  wire [31:0] x429_sum_1_io_result; // @[Math.scala 150:24:@28642.4]
  wire  x432_sum_1_clock; // @[Math.scala 150:24:@28680.4]
  wire  x432_sum_1_reset; // @[Math.scala 150:24:@28680.4]
  wire [31:0] x432_sum_1_io_a; // @[Math.scala 150:24:@28680.4]
  wire [31:0] x432_sum_1_io_b; // @[Math.scala 150:24:@28680.4]
  wire  x432_sum_1_io_flow; // @[Math.scala 150:24:@28680.4]
  wire [31:0] x432_sum_1_io_result; // @[Math.scala 150:24:@28680.4]
  wire  x435_sum_1_clock; // @[Math.scala 150:24:@28718.4]
  wire  x435_sum_1_reset; // @[Math.scala 150:24:@28718.4]
  wire [31:0] x435_sum_1_io_a; // @[Math.scala 150:24:@28718.4]
  wire [31:0] x435_sum_1_io_b; // @[Math.scala 150:24:@28718.4]
  wire  x435_sum_1_io_flow; // @[Math.scala 150:24:@28718.4]
  wire [31:0] x435_sum_1_io_result; // @[Math.scala 150:24:@28718.4]
  wire  x438_sum_1_clock; // @[Math.scala 150:24:@28756.4]
  wire  x438_sum_1_reset; // @[Math.scala 150:24:@28756.4]
  wire [31:0] x438_sum_1_io_a; // @[Math.scala 150:24:@28756.4]
  wire [31:0] x438_sum_1_io_b; // @[Math.scala 150:24:@28756.4]
  wire  x438_sum_1_io_flow; // @[Math.scala 150:24:@28756.4]
  wire [31:0] x438_sum_1_io_result; // @[Math.scala 150:24:@28756.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@28771.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@28771.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@28771.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@28771.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@28771.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@28785.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@28785.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@28785.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@28785.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@28785.4]
  wire  x441_sub_1_clock; // @[Math.scala 191:24:@28796.4]
  wire  x441_sub_1_reset; // @[Math.scala 191:24:@28796.4]
  wire [31:0] x441_sub_1_io_a; // @[Math.scala 191:24:@28796.4]
  wire [31:0] x441_sub_1_io_b; // @[Math.scala 191:24:@28796.4]
  wire  x441_sub_1_io_flow; // @[Math.scala 191:24:@28796.4]
  wire [31:0] x441_sub_1_io_result; // @[Math.scala 191:24:@28796.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@28806.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@28806.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@28806.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@28806.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@28806.4]
  wire  x250_div_1_clock; // @[Math.scala 327:24:@28820.4]
  wire [31:0] x250_div_1_io_a; // @[Math.scala 327:24:@28820.4]
  wire  x250_div_1_io_flow; // @[Math.scala 327:24:@28820.4]
  wire [31:0] x250_div_1_io_result; // @[Math.scala 327:24:@28820.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@28830.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@28830.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@28830.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@28830.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@28830.4]
  wire  x251_sum_1_clock; // @[Math.scala 150:24:@28839.4]
  wire  x251_sum_1_reset; // @[Math.scala 150:24:@28839.4]
  wire [31:0] x251_sum_1_io_a; // @[Math.scala 150:24:@28839.4]
  wire [31:0] x251_sum_1_io_b; // @[Math.scala 150:24:@28839.4]
  wire  x251_sum_1_io_flow; // @[Math.scala 150:24:@28839.4]
  wire [31:0] x251_sum_1_io_result; // @[Math.scala 150:24:@28839.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@28849.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@28849.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@28849.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@28849.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@28849.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@28858.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@28858.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@28858.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@28858.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@28858.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@28870.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@28870.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@28870.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@28870.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@28870.4]
  wire  x254_rdcol_1_clock; // @[Math.scala 191:24:@28893.4]
  wire  x254_rdcol_1_reset; // @[Math.scala 191:24:@28893.4]
  wire [31:0] x254_rdcol_1_io_a; // @[Math.scala 191:24:@28893.4]
  wire [31:0] x254_rdcol_1_io_b; // @[Math.scala 191:24:@28893.4]
  wire  x254_rdcol_1_io_flow; // @[Math.scala 191:24:@28893.4]
  wire [31:0] x254_rdcol_1_io_result; // @[Math.scala 191:24:@28893.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@28908.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@28908.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@28908.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@28908.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@28908.4]
  wire  x445_sum_1_clock; // @[Math.scala 150:24:@28953.4]
  wire  x445_sum_1_reset; // @[Math.scala 150:24:@28953.4]
  wire [31:0] x445_sum_1_io_a; // @[Math.scala 150:24:@28953.4]
  wire [31:0] x445_sum_1_io_b; // @[Math.scala 150:24:@28953.4]
  wire  x445_sum_1_io_flow; // @[Math.scala 150:24:@28953.4]
  wire [31:0] x445_sum_1_io_result; // @[Math.scala 150:24:@28953.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@28976.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@28976.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@28976.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@28976.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@28976.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@28994.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@28994.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@28994.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@28994.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@28994.4]
  wire  x448_sum_1_clock; // @[Math.scala 150:24:@29007.4]
  wire  x448_sum_1_reset; // @[Math.scala 150:24:@29007.4]
  wire [31:0] x448_sum_1_io_a; // @[Math.scala 150:24:@29007.4]
  wire [31:0] x448_sum_1_io_b; // @[Math.scala 150:24:@29007.4]
  wire  x448_sum_1_io_flow; // @[Math.scala 150:24:@29007.4]
  wire [31:0] x448_sum_1_io_result; // @[Math.scala 150:24:@29007.4]
  wire  x451_sum_1_clock; // @[Math.scala 150:24:@29045.4]
  wire  x451_sum_1_reset; // @[Math.scala 150:24:@29045.4]
  wire [31:0] x451_sum_1_io_a; // @[Math.scala 150:24:@29045.4]
  wire [31:0] x451_sum_1_io_b; // @[Math.scala 150:24:@29045.4]
  wire  x451_sum_1_io_flow; // @[Math.scala 150:24:@29045.4]
  wire [31:0] x451_sum_1_io_result; // @[Math.scala 150:24:@29045.4]
  wire  x454_sum_1_clock; // @[Math.scala 150:24:@29083.4]
  wire  x454_sum_1_reset; // @[Math.scala 150:24:@29083.4]
  wire [31:0] x454_sum_1_io_a; // @[Math.scala 150:24:@29083.4]
  wire [31:0] x454_sum_1_io_b; // @[Math.scala 150:24:@29083.4]
  wire  x454_sum_1_io_flow; // @[Math.scala 150:24:@29083.4]
  wire [31:0] x454_sum_1_io_result; // @[Math.scala 150:24:@29083.4]
  wire  x457_sum_1_clock; // @[Math.scala 150:24:@29121.4]
  wire  x457_sum_1_reset; // @[Math.scala 150:24:@29121.4]
  wire [31:0] x457_sum_1_io_a; // @[Math.scala 150:24:@29121.4]
  wire [31:0] x457_sum_1_io_b; // @[Math.scala 150:24:@29121.4]
  wire  x457_sum_1_io_flow; // @[Math.scala 150:24:@29121.4]
  wire [31:0] x457_sum_1_io_result; // @[Math.scala 150:24:@29121.4]
  wire  x460_sum_1_clock; // @[Math.scala 150:24:@29159.4]
  wire  x460_sum_1_reset; // @[Math.scala 150:24:@29159.4]
  wire [31:0] x460_sum_1_io_a; // @[Math.scala 150:24:@29159.4]
  wire [31:0] x460_sum_1_io_b; // @[Math.scala 150:24:@29159.4]
  wire  x460_sum_1_io_flow; // @[Math.scala 150:24:@29159.4]
  wire [31:0] x460_sum_1_io_result; // @[Math.scala 150:24:@29159.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@29174.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@29174.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@29174.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@29174.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@29174.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@29188.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@29188.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@29188.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@29188.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@29188.4]
  wire  x463_sub_1_clock; // @[Math.scala 191:24:@29199.4]
  wire  x463_sub_1_reset; // @[Math.scala 191:24:@29199.4]
  wire [31:0] x463_sub_1_io_a; // @[Math.scala 191:24:@29199.4]
  wire [31:0] x463_sub_1_io_b; // @[Math.scala 191:24:@29199.4]
  wire  x463_sub_1_io_flow; // @[Math.scala 191:24:@29199.4]
  wire [31:0] x463_sub_1_io_result; // @[Math.scala 191:24:@29199.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@29209.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@29209.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@29209.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@29209.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@29209.4]
  wire  x259_div_1_clock; // @[Math.scala 327:24:@29223.4]
  wire [31:0] x259_div_1_io_a; // @[Math.scala 327:24:@29223.4]
  wire  x259_div_1_io_flow; // @[Math.scala 327:24:@29223.4]
  wire [31:0] x259_div_1_io_result; // @[Math.scala 327:24:@29223.4]
  wire  x260_sum_1_clock; // @[Math.scala 150:24:@29233.4]
  wire  x260_sum_1_reset; // @[Math.scala 150:24:@29233.4]
  wire [31:0] x260_sum_1_io_a; // @[Math.scala 150:24:@29233.4]
  wire [31:0] x260_sum_1_io_b; // @[Math.scala 150:24:@29233.4]
  wire  x260_sum_1_io_flow; // @[Math.scala 150:24:@29233.4]
  wire [31:0] x260_sum_1_io_result; // @[Math.scala 150:24:@29233.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@29243.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@29252.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@29252.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@29252.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@29264.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@29264.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@29264.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@29264.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@29264.4]
  wire  x263_rdrow_1_clock; // @[Math.scala 191:24:@29287.4]
  wire  x263_rdrow_1_reset; // @[Math.scala 191:24:@29287.4]
  wire [31:0] x263_rdrow_1_io_a; // @[Math.scala 191:24:@29287.4]
  wire [31:0] x263_rdrow_1_io_b; // @[Math.scala 191:24:@29287.4]
  wire  x263_rdrow_1_io_flow; // @[Math.scala 191:24:@29287.4]
  wire [31:0] x263_rdrow_1_io_result; // @[Math.scala 191:24:@29287.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@29313.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@29313.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@29313.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@29313.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@29313.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@29322.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@29322.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@29322.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@29322.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@29322.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@29344.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@29344.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@29344.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@29344.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@29344.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@29370.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@29370.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@29370.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@29370.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@29370.4]
  wire  x469_sum_1_clock; // @[Math.scala 150:24:@29391.4]
  wire  x469_sum_1_reset; // @[Math.scala 150:24:@29391.4]
  wire [31:0] x469_sum_1_io_a; // @[Math.scala 150:24:@29391.4]
  wire [31:0] x469_sum_1_io_b; // @[Math.scala 150:24:@29391.4]
  wire  x469_sum_1_io_flow; // @[Math.scala 150:24:@29391.4]
  wire [31:0] x469_sum_1_io_result; // @[Math.scala 150:24:@29391.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@29401.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@29401.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@29401.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@29401.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@29401.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@29410.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@29410.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@29410.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@29410.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@29410.4]
  wire  x271_sum_1_clock; // @[Math.scala 150:24:@29419.4]
  wire  x271_sum_1_reset; // @[Math.scala 150:24:@29419.4]
  wire [31:0] x271_sum_1_io_a; // @[Math.scala 150:24:@29419.4]
  wire [31:0] x271_sum_1_io_b; // @[Math.scala 150:24:@29419.4]
  wire  x271_sum_1_io_flow; // @[Math.scala 150:24:@29419.4]
  wire [31:0] x271_sum_1_io_result; // @[Math.scala 150:24:@29419.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@29429.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@29429.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@29429.4]
  wire [31:0] RetimeWrapper_50_io_in; // @[package.scala 93:22:@29429.4]
  wire [31:0] RetimeWrapper_50_io_out; // @[package.scala 93:22:@29429.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@29438.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@29438.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@29438.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@29438.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@29438.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@29447.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@29447.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@29447.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@29447.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@29447.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@29459.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@29459.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@29459.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@29459.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@29459.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@29486.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@29486.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@29486.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@29486.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@29486.4]
  wire  x276_sum_1_clock; // @[Math.scala 150:24:@29497.4]
  wire  x276_sum_1_reset; // @[Math.scala 150:24:@29497.4]
  wire [31:0] x276_sum_1_io_a; // @[Math.scala 150:24:@29497.4]
  wire [31:0] x276_sum_1_io_b; // @[Math.scala 150:24:@29497.4]
  wire  x276_sum_1_io_flow; // @[Math.scala 150:24:@29497.4]
  wire [31:0] x276_sum_1_io_result; // @[Math.scala 150:24:@29497.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@29507.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@29507.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@29507.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@29507.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@29507.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@29519.4]
  wire  x281_sum_1_clock; // @[Math.scala 150:24:@29546.4]
  wire  x281_sum_1_reset; // @[Math.scala 150:24:@29546.4]
  wire [31:0] x281_sum_1_io_a; // @[Math.scala 150:24:@29546.4]
  wire [31:0] x281_sum_1_io_b; // @[Math.scala 150:24:@29546.4]
  wire  x281_sum_1_io_flow; // @[Math.scala 150:24:@29546.4]
  wire [31:0] x281_sum_1_io_result; // @[Math.scala 150:24:@29546.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@29556.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@29556.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@29556.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@29556.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@29556.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@29568.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@29568.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@29568.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@29568.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@29568.4]
  wire  x284_rdrow_1_clock; // @[Math.scala 191:24:@29591.4]
  wire  x284_rdrow_1_reset; // @[Math.scala 191:24:@29591.4]
  wire [31:0] x284_rdrow_1_io_a; // @[Math.scala 191:24:@29591.4]
  wire [31:0] x284_rdrow_1_io_b; // @[Math.scala 191:24:@29591.4]
  wire  x284_rdrow_1_io_flow; // @[Math.scala 191:24:@29591.4]
  wire [31:0] x284_rdrow_1_io_result; // @[Math.scala 191:24:@29591.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@29617.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@29617.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@29617.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@29617.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@29617.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@29639.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@29639.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@29639.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@29639.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@29639.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@29665.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@29665.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@29665.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@29665.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@29665.4]
  wire  x474_sum_1_clock; // @[Math.scala 150:24:@29686.4]
  wire  x474_sum_1_reset; // @[Math.scala 150:24:@29686.4]
  wire [31:0] x474_sum_1_io_a; // @[Math.scala 150:24:@29686.4]
  wire [31:0] x474_sum_1_io_b; // @[Math.scala 150:24:@29686.4]
  wire  x474_sum_1_io_flow; // @[Math.scala 150:24:@29686.4]
  wire [31:0] x474_sum_1_io_result; // @[Math.scala 150:24:@29686.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@29696.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@29696.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@29696.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@29696.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@29696.4]
  wire  x292_sum_1_clock; // @[Math.scala 150:24:@29705.4]
  wire  x292_sum_1_reset; // @[Math.scala 150:24:@29705.4]
  wire [31:0] x292_sum_1_io_a; // @[Math.scala 150:24:@29705.4]
  wire [31:0] x292_sum_1_io_b; // @[Math.scala 150:24:@29705.4]
  wire  x292_sum_1_io_flow; // @[Math.scala 150:24:@29705.4]
  wire [31:0] x292_sum_1_io_result; // @[Math.scala 150:24:@29705.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@29715.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@29715.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@29715.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@29715.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@29715.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@29724.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@29724.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@29724.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@29724.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@29724.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@29733.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@29733.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@29733.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@29733.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@29733.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@29745.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@29745.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@29745.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@29745.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@29745.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@29772.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@29772.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@29772.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@29772.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@29772.4]
  wire  x297_sum_1_clock; // @[Math.scala 150:24:@29781.4]
  wire  x297_sum_1_reset; // @[Math.scala 150:24:@29781.4]
  wire [31:0] x297_sum_1_io_a; // @[Math.scala 150:24:@29781.4]
  wire [31:0] x297_sum_1_io_b; // @[Math.scala 150:24:@29781.4]
  wire  x297_sum_1_io_flow; // @[Math.scala 150:24:@29781.4]
  wire [31:0] x297_sum_1_io_result; // @[Math.scala 150:24:@29781.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@29791.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@29791.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@29791.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@29791.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@29791.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@29803.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@29803.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@29803.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@29803.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@29803.4]
  wire  x302_sum_1_clock; // @[Math.scala 150:24:@29830.4]
  wire  x302_sum_1_reset; // @[Math.scala 150:24:@29830.4]
  wire [31:0] x302_sum_1_io_a; // @[Math.scala 150:24:@29830.4]
  wire [31:0] x302_sum_1_io_b; // @[Math.scala 150:24:@29830.4]
  wire  x302_sum_1_io_flow; // @[Math.scala 150:24:@29830.4]
  wire [31:0] x302_sum_1_io_result; // @[Math.scala 150:24:@29830.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@29840.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@29840.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@29840.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@29840.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@29840.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@29852.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@29852.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@29852.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@29852.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@29852.4]
  wire  x305_1_clock; // @[Math.scala 262:24:@29875.4]
  wire [31:0] x305_1_io_a; // @[Math.scala 262:24:@29875.4]
  wire [31:0] x305_1_io_b; // @[Math.scala 262:24:@29875.4]
  wire  x305_1_io_flow; // @[Math.scala 262:24:@29875.4]
  wire [31:0] x305_1_io_result; // @[Math.scala 262:24:@29875.4]
  wire  x306_1_clock; // @[Math.scala 262:24:@29887.4]
  wire [31:0] x306_1_io_a; // @[Math.scala 262:24:@29887.4]
  wire [31:0] x306_1_io_b; // @[Math.scala 262:24:@29887.4]
  wire  x306_1_io_flow; // @[Math.scala 262:24:@29887.4]
  wire [31:0] x306_1_io_result; // @[Math.scala 262:24:@29887.4]
  wire  x307_1_clock; // @[Math.scala 262:24:@29899.4]
  wire [31:0] x307_1_io_a; // @[Math.scala 262:24:@29899.4]
  wire [31:0] x307_1_io_b; // @[Math.scala 262:24:@29899.4]
  wire  x307_1_io_flow; // @[Math.scala 262:24:@29899.4]
  wire [31:0] x307_1_io_result; // @[Math.scala 262:24:@29899.4]
  wire  x308_1_clock; // @[Math.scala 262:24:@29911.4]
  wire [31:0] x308_1_io_a; // @[Math.scala 262:24:@29911.4]
  wire [31:0] x308_1_io_b; // @[Math.scala 262:24:@29911.4]
  wire  x308_1_io_flow; // @[Math.scala 262:24:@29911.4]
  wire [31:0] x308_1_io_result; // @[Math.scala 262:24:@29911.4]
  wire  x309_1_clock; // @[Math.scala 262:24:@29923.4]
  wire [31:0] x309_1_io_a; // @[Math.scala 262:24:@29923.4]
  wire [31:0] x309_1_io_b; // @[Math.scala 262:24:@29923.4]
  wire  x309_1_io_flow; // @[Math.scala 262:24:@29923.4]
  wire [31:0] x309_1_io_result; // @[Math.scala 262:24:@29923.4]
  wire  x310_1_clock; // @[Math.scala 262:24:@29937.4]
  wire [31:0] x310_1_io_a; // @[Math.scala 262:24:@29937.4]
  wire [31:0] x310_1_io_b; // @[Math.scala 262:24:@29937.4]
  wire  x310_1_io_flow; // @[Math.scala 262:24:@29937.4]
  wire [31:0] x310_1_io_result; // @[Math.scala 262:24:@29937.4]
  wire  x311_1_clock; // @[Math.scala 262:24:@29949.4]
  wire [31:0] x311_1_io_a; // @[Math.scala 262:24:@29949.4]
  wire [31:0] x311_1_io_b; // @[Math.scala 262:24:@29949.4]
  wire  x311_1_io_flow; // @[Math.scala 262:24:@29949.4]
  wire [31:0] x311_1_io_result; // @[Math.scala 262:24:@29949.4]
  wire  x312_1_clock; // @[Math.scala 262:24:@29961.4]
  wire [31:0] x312_1_io_a; // @[Math.scala 262:24:@29961.4]
  wire [31:0] x312_1_io_b; // @[Math.scala 262:24:@29961.4]
  wire  x312_1_io_flow; // @[Math.scala 262:24:@29961.4]
  wire [31:0] x312_1_io_result; // @[Math.scala 262:24:@29961.4]
  wire  x313_1_clock; // @[Math.scala 262:24:@29973.4]
  wire [31:0] x313_1_io_a; // @[Math.scala 262:24:@29973.4]
  wire [31:0] x313_1_io_b; // @[Math.scala 262:24:@29973.4]
  wire  x313_1_io_flow; // @[Math.scala 262:24:@29973.4]
  wire [31:0] x313_1_io_result; // @[Math.scala 262:24:@29973.4]
  wire  x314_x13_1_clock; // @[Math.scala 150:24:@29983.4]
  wire  x314_x13_1_reset; // @[Math.scala 150:24:@29983.4]
  wire [31:0] x314_x13_1_io_a; // @[Math.scala 150:24:@29983.4]
  wire [31:0] x314_x13_1_io_b; // @[Math.scala 150:24:@29983.4]
  wire  x314_x13_1_io_flow; // @[Math.scala 150:24:@29983.4]
  wire [31:0] x314_x13_1_io_result; // @[Math.scala 150:24:@29983.4]
  wire  x315_x14_1_clock; // @[Math.scala 150:24:@29993.4]
  wire  x315_x14_1_reset; // @[Math.scala 150:24:@29993.4]
  wire [31:0] x315_x14_1_io_a; // @[Math.scala 150:24:@29993.4]
  wire [31:0] x315_x14_1_io_b; // @[Math.scala 150:24:@29993.4]
  wire  x315_x14_1_io_flow; // @[Math.scala 150:24:@29993.4]
  wire [31:0] x315_x14_1_io_result; // @[Math.scala 150:24:@29993.4]
  wire  x316_x13_1_clock; // @[Math.scala 150:24:@30003.4]
  wire  x316_x13_1_reset; // @[Math.scala 150:24:@30003.4]
  wire [31:0] x316_x13_1_io_a; // @[Math.scala 150:24:@30003.4]
  wire [31:0] x316_x13_1_io_b; // @[Math.scala 150:24:@30003.4]
  wire  x316_x13_1_io_flow; // @[Math.scala 150:24:@30003.4]
  wire [31:0] x316_x13_1_io_result; // @[Math.scala 150:24:@30003.4]
  wire  x317_x14_1_clock; // @[Math.scala 150:24:@30013.4]
  wire  x317_x14_1_reset; // @[Math.scala 150:24:@30013.4]
  wire [31:0] x317_x14_1_io_a; // @[Math.scala 150:24:@30013.4]
  wire [31:0] x317_x14_1_io_b; // @[Math.scala 150:24:@30013.4]
  wire  x317_x14_1_io_flow; // @[Math.scala 150:24:@30013.4]
  wire [31:0] x317_x14_1_io_result; // @[Math.scala 150:24:@30013.4]
  wire  x318_x13_1_clock; // @[Math.scala 150:24:@30023.4]
  wire  x318_x13_1_reset; // @[Math.scala 150:24:@30023.4]
  wire [31:0] x318_x13_1_io_a; // @[Math.scala 150:24:@30023.4]
  wire [31:0] x318_x13_1_io_b; // @[Math.scala 150:24:@30023.4]
  wire  x318_x13_1_io_flow; // @[Math.scala 150:24:@30023.4]
  wire [31:0] x318_x13_1_io_result; // @[Math.scala 150:24:@30023.4]
  wire  x319_x14_1_clock; // @[Math.scala 150:24:@30033.4]
  wire  x319_x14_1_reset; // @[Math.scala 150:24:@30033.4]
  wire [31:0] x319_x14_1_io_a; // @[Math.scala 150:24:@30033.4]
  wire [31:0] x319_x14_1_io_b; // @[Math.scala 150:24:@30033.4]
  wire  x319_x14_1_io_flow; // @[Math.scala 150:24:@30033.4]
  wire [31:0] x319_x14_1_io_result; // @[Math.scala 150:24:@30033.4]
  wire  x320_x13_1_clock; // @[Math.scala 150:24:@30043.4]
  wire  x320_x13_1_reset; // @[Math.scala 150:24:@30043.4]
  wire [31:0] x320_x13_1_io_a; // @[Math.scala 150:24:@30043.4]
  wire [31:0] x320_x13_1_io_b; // @[Math.scala 150:24:@30043.4]
  wire  x320_x13_1_io_flow; // @[Math.scala 150:24:@30043.4]
  wire [31:0] x320_x13_1_io_result; // @[Math.scala 150:24:@30043.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@30053.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@30053.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@30053.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@30053.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@30053.4]
  wire  x321_sum_1_clock; // @[Math.scala 150:24:@30062.4]
  wire  x321_sum_1_reset; // @[Math.scala 150:24:@30062.4]
  wire [31:0] x321_sum_1_io_a; // @[Math.scala 150:24:@30062.4]
  wire [31:0] x321_sum_1_io_b; // @[Math.scala 150:24:@30062.4]
  wire  x321_sum_1_io_flow; // @[Math.scala 150:24:@30062.4]
  wire [31:0] x321_sum_1_io_result; // @[Math.scala 150:24:@30062.4]
  wire [31:0] x322_1_io_b; // @[Math.scala 720:24:@30072.4]
  wire [31:0] x322_1_io_result; // @[Math.scala 720:24:@30072.4]
  wire  x323_mul_1_clock; // @[Math.scala 262:24:@30083.4]
  wire [31:0] x323_mul_1_io_a; // @[Math.scala 262:24:@30083.4]
  wire [31:0] x323_mul_1_io_b; // @[Math.scala 262:24:@30083.4]
  wire  x323_mul_1_io_flow; // @[Math.scala 262:24:@30083.4]
  wire [31:0] x323_mul_1_io_result; // @[Math.scala 262:24:@30083.4]
  wire [31:0] x324_1_io_b; // @[Math.scala 720:24:@30093.4]
  wire [31:0] x324_1_io_result; // @[Math.scala 720:24:@30093.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@30102.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@30102.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@30102.4]
  wire [31:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@30102.4]
  wire [31:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@30102.4]
  wire  x325_sub_1_clock; // @[Math.scala 191:24:@30111.4]
  wire  x325_sub_1_reset; // @[Math.scala 191:24:@30111.4]
  wire [31:0] x325_sub_1_io_a; // @[Math.scala 191:24:@30111.4]
  wire [31:0] x325_sub_1_io_b; // @[Math.scala 191:24:@30111.4]
  wire  x325_sub_1_io_flow; // @[Math.scala 191:24:@30111.4]
  wire [31:0] x325_sub_1_io_result; // @[Math.scala 191:24:@30111.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@30124.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@30124.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@30124.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@30124.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@30124.4]
  wire  x327_sub_1_clock; // @[Math.scala 191:24:@30133.4]
  wire  x327_sub_1_reset; // @[Math.scala 191:24:@30133.4]
  wire [31:0] x327_sub_1_io_a; // @[Math.scala 191:24:@30133.4]
  wire [31:0] x327_sub_1_io_b; // @[Math.scala 191:24:@30133.4]
  wire  x327_sub_1_io_flow; // @[Math.scala 191:24:@30133.4]
  wire [31:0] x327_sub_1_io_result; // @[Math.scala 191:24:@30133.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@30146.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@30146.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@30146.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@30146.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@30146.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@30158.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@30158.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@30158.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@30158.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@30158.4]
  wire [31:0] x331_1_io_b; // @[Math.scala 720:24:@30172.4]
  wire [31:0] x331_1_io_result; // @[Math.scala 720:24:@30172.4]
  wire  x332_mul_1_clock; // @[Math.scala 262:24:@30183.4]
  wire [31:0] x332_mul_1_io_a; // @[Math.scala 262:24:@30183.4]
  wire [31:0] x332_mul_1_io_b; // @[Math.scala 262:24:@30183.4]
  wire  x332_mul_1_io_flow; // @[Math.scala 262:24:@30183.4]
  wire [31:0] x332_mul_1_io_result; // @[Math.scala 262:24:@30183.4]
  wire [31:0] x333_1_io_b; // @[Math.scala 720:24:@30193.4]
  wire [31:0] x333_1_io_result; // @[Math.scala 720:24:@30193.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@30202.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@30202.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@30202.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@30202.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@30202.4]
  wire  x334_sum_1_clock; // @[Math.scala 150:24:@30211.4]
  wire  x334_sum_1_reset; // @[Math.scala 150:24:@30211.4]
  wire [31:0] x334_sum_1_io_a; // @[Math.scala 150:24:@30211.4]
  wire [31:0] x334_sum_1_io_b; // @[Math.scala 150:24:@30211.4]
  wire  x334_sum_1_io_flow; // @[Math.scala 150:24:@30211.4]
  wire [31:0] x334_sum_1_io_result; // @[Math.scala 150:24:@30211.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@30225.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@30225.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@30225.4]
  wire [31:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@30225.4]
  wire [31:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@30225.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@30234.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@30234.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@30234.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@30234.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@30234.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@30252.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@30252.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@30252.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@30252.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@30252.4]
  wire  b223; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 62:18:@27791.4]
  wire  b224; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 63:18:@27792.4]
  wire  _T_205; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 67:30:@27794.4]
  wire  _T_206; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 67:37:@27795.4]
  wire  _T_210; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 69:76:@27800.4]
  wire  _T_211; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 69:62:@27801.4]
  wire  _T_213; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 69:101:@27802.4]
  wire [31:0] b221_number; // @[Math.scala 723:22:@27776.4 Math.scala 724:14:@27777.4]
  wire [31:0] _T_241; // @[Math.scala 406:49:@27892.4]
  wire [31:0] _T_243; // @[Math.scala 406:56:@27894.4]
  wire [31:0] _T_244; // @[Math.scala 406:56:@27895.4]
  wire [31:0] x394_number; // @[implicits.scala 133:21:@27896.4]
  wire [31:0] _T_254; // @[Math.scala 406:49:@27905.4]
  wire [31:0] _T_256; // @[Math.scala 406:56:@27907.4]
  wire [31:0] _T_257; // @[Math.scala 406:56:@27908.4]
  wire [31:0] b222_number; // @[Math.scala 723:22:@27788.4 Math.scala 724:14:@27789.4]
  wire  _T_261; // @[FixedPoint.scala 50:25:@27914.4]
  wire [15:0] _T_265; // @[Bitwise.scala 72:12:@27916.4]
  wire [15:0] _T_266; // @[FixedPoint.scala 18:52:@27917.4]
  wire  _T_272; // @[Math.scala 451:55:@27919.4]
  wire [15:0] _T_273; // @[FixedPoint.scala 18:52:@27920.4]
  wire  _T_279; // @[Math.scala 451:110:@27922.4]
  wire  _T_280; // @[Math.scala 451:94:@27923.4]
  wire [31:0] _T_282; // @[Cat.scala 30:58:@27925.4]
  wire [31:0] _T_292; // @[Math.scala 406:49:@27933.4]
  wire [31:0] _T_294; // @[Math.scala 406:56:@27935.4]
  wire [31:0] _T_295; // @[Math.scala 406:56:@27936.4]
  wire [31:0] x398_sum_number; // @[Math.scala 154:22:@27947.4 Math.scala 155:14:@27948.4]
  wire  _T_302; // @[FixedPoint.scala 50:25:@27952.4]
  wire [7:0] _T_306; // @[Bitwise.scala 72:12:@27954.4]
  wire [23:0] _T_307; // @[FixedPoint.scala 18:52:@27955.4]
  wire  _T_313; // @[Math.scala 451:55:@27957.4]
  wire [7:0] _T_314; // @[FixedPoint.scala 18:52:@27958.4]
  wire  _T_320; // @[Math.scala 451:110:@27960.4]
  wire  _T_321; // @[Math.scala 451:94:@27961.4]
  wire [31:0] _T_323; // @[Cat.scala 30:58:@27963.4]
  wire [31:0] _T_333; // @[Math.scala 406:49:@27971.4]
  wire [31:0] _T_335; // @[Math.scala 406:56:@27973.4]
  wire [31:0] _T_336; // @[Math.scala 406:56:@27974.4]
  wire [31:0] x401_sum_number; // @[Math.scala 154:22:@27985.4 Math.scala 155:14:@27986.4]
  wire  _T_343; // @[FixedPoint.scala 50:25:@27990.4]
  wire [3:0] _T_347; // @[Bitwise.scala 72:12:@27992.4]
  wire [27:0] _T_348; // @[FixedPoint.scala 18:52:@27993.4]
  wire  _T_354; // @[Math.scala 451:55:@27995.4]
  wire [3:0] _T_355; // @[FixedPoint.scala 18:52:@27996.4]
  wire  _T_361; // @[Math.scala 451:110:@27998.4]
  wire  _T_362; // @[Math.scala 451:94:@27999.4]
  wire [31:0] _T_364; // @[Cat.scala 30:58:@28001.4]
  wire [31:0] _T_374; // @[Math.scala 406:49:@28009.4]
  wire [31:0] _T_376; // @[Math.scala 406:56:@28011.4]
  wire [31:0] _T_377; // @[Math.scala 406:56:@28012.4]
  wire [31:0] x404_sum_number; // @[Math.scala 154:22:@28023.4 Math.scala 155:14:@28024.4]
  wire  _T_384; // @[FixedPoint.scala 50:25:@28028.4]
  wire [1:0] _T_388; // @[Bitwise.scala 72:12:@28030.4]
  wire [29:0] _T_389; // @[FixedPoint.scala 18:52:@28031.4]
  wire  _T_395; // @[Math.scala 451:55:@28033.4]
  wire [1:0] _T_396; // @[FixedPoint.scala 18:52:@28034.4]
  wire  _T_402; // @[Math.scala 451:110:@28036.4]
  wire  _T_403; // @[Math.scala 451:94:@28037.4]
  wire [31:0] _T_405; // @[Cat.scala 30:58:@28039.4]
  wire [31:0] _T_415; // @[Math.scala 406:49:@28047.4]
  wire [31:0] _T_417; // @[Math.scala 406:56:@28049.4]
  wire [31:0] _T_418; // @[Math.scala 406:56:@28050.4]
  wire [31:0] x407_sum_number; // @[Math.scala 154:22:@28061.4 Math.scala 155:14:@28062.4]
  wire  _T_425; // @[FixedPoint.scala 50:25:@28066.4]
  wire [1:0] _T_429; // @[Bitwise.scala 72:12:@28068.4]
  wire [29:0] _T_430; // @[FixedPoint.scala 18:52:@28069.4]
  wire  _T_436; // @[Math.scala 451:55:@28071.4]
  wire [1:0] _T_437; // @[FixedPoint.scala 18:52:@28072.4]
  wire  _T_443; // @[Math.scala 451:110:@28074.4]
  wire  _T_444; // @[Math.scala 451:94:@28075.4]
  wire [31:0] _T_448; // @[package.scala 96:25:@28083.4 package.scala 96:25:@28084.4]
  wire [31:0] _T_458; // @[Math.scala 406:49:@28092.4]
  wire [31:0] _T_460; // @[Math.scala 406:56:@28094.4]
  wire [31:0] _T_461; // @[Math.scala 406:56:@28095.4]
  wire [31:0] _T_465; // @[package.scala 96:25:@28103.4]
  wire [31:0] x410_sum_number; // @[Math.scala 154:22:@28115.4 Math.scala 155:14:@28116.4]
  wire  _T_472; // @[FixedPoint.scala 50:25:@28120.4]
  wire [1:0] _T_476; // @[Bitwise.scala 72:12:@28122.4]
  wire [29:0] _T_477; // @[FixedPoint.scala 18:52:@28123.4]
  wire  _T_483; // @[Math.scala 451:55:@28125.4]
  wire [1:0] _T_484; // @[FixedPoint.scala 18:52:@28126.4]
  wire  _T_490; // @[Math.scala 451:110:@28128.4]
  wire  _T_491; // @[Math.scala 451:94:@28129.4]
  wire [31:0] _T_493; // @[Cat.scala 30:58:@28131.4]
  wire [31:0] _T_503; // @[Math.scala 406:49:@28139.4]
  wire [31:0] _T_505; // @[Math.scala 406:56:@28141.4]
  wire [31:0] _T_506; // @[Math.scala 406:56:@28142.4]
  wire [31:0] x413_sum_number; // @[Math.scala 154:22:@28153.4 Math.scala 155:14:@28154.4]
  wire [31:0] _T_516; // @[Math.scala 476:37:@28159.4]
  wire  x482_x414_D1; // @[package.scala 96:25:@28197.4 package.scala 96:25:@28198.4]
  wire [31:0] x483_x413_sum_D1_number; // @[package.scala 96:25:@28206.4 package.scala 96:25:@28207.4]
  wire [31:0] x416_sub_number; // @[Math.scala 195:22:@28179.4 Math.scala 196:14:@28180.4]
  wire  _T_547; // @[FixedPoint.scala 50:25:@28214.4]
  wire [1:0] _T_551; // @[Bitwise.scala 72:12:@28216.4]
  wire [29:0] _T_552; // @[FixedPoint.scala 18:52:@28217.4]
  wire  _T_558; // @[Math.scala 451:55:@28219.4]
  wire [1:0] _T_559; // @[FixedPoint.scala 18:52:@28220.4]
  wire  _T_565; // @[Math.scala 451:110:@28222.4]
  wire  _T_566; // @[Math.scala 451:94:@28223.4]
  wire [31:0] _T_568; // @[Cat.scala 30:58:@28225.4]
  wire [31:0] x233_1_number; // @[Math.scala 454:20:@28226.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@28231.4]
  wire [40:0] _T_573; // @[Math.scala 461:32:@28231.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@28236.4]
  wire [38:0] _T_576; // @[Math.scala 461:32:@28236.4]
  wire  _T_609; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:101:@28325.4]
  wire  _T_613; // @[package.scala 96:25:@28333.4 package.scala 96:25:@28334.4]
  wire  _T_615; // @[implicits.scala 55:10:@28335.4]
  wire  _T_616; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:118:@28336.4]
  wire  _T_618; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:207:@28338.4]
  wire  _T_619; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:226:@28339.4]
  wire  x488_b223_D21; // @[package.scala 96:25:@28313.4 package.scala 96:25:@28314.4]
  wire  _T_620; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:252:@28340.4]
  wire  x486_b224_D21; // @[package.scala 96:25:@28295.4 package.scala 96:25:@28296.4]
  wire [31:0] x490_b221_D23_number; // @[package.scala 96:25:@28354.4 package.scala 96:25:@28355.4]
  wire [31:0] _T_630; // @[Math.scala 476:37:@28360.4]
  wire [31:0] x491_b222_D23_number; // @[package.scala 96:25:@28377.4 package.scala 96:25:@28378.4]
  wire [31:0] _T_645; // @[Math.scala 476:37:@28385.4]
  wire  x239; // @[package.scala 96:25:@28368.4 package.scala 96:25:@28369.4]
  wire  x240; // @[package.scala 96:25:@28393.4 package.scala 96:25:@28394.4]
  wire  x241; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 182:59:@28397.4]
  wire  _T_683; // @[package.scala 96:25:@28465.4 package.scala 96:25:@28466.4]
  wire  _T_685; // @[implicits.scala 55:10:@28467.4]
  wire  _T_686; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 201:194:@28468.4]
  wire  x496_x242_D21; // @[package.scala 96:25:@28444.4 package.scala 96:25:@28445.4]
  wire  _T_687; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 201:283:@28469.4]
  wire  x495_b223_D45; // @[package.scala 96:25:@28435.4 package.scala 96:25:@28436.4]
  wire  _T_688; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 201:291:@28470.4]
  wire  x493_b224_D45; // @[package.scala 96:25:@28417.4 package.scala 96:25:@28418.4]
  wire [31:0] x245_rdcol_number; // @[Math.scala 195:22:@28489.4 Math.scala 196:14:@28490.4]
  wire [31:0] _T_703; // @[Math.scala 476:37:@28495.4]
  wire  x498_x239_D1; // @[package.scala 96:25:@28512.4 package.scala 96:25:@28513.4]
  wire  x246; // @[package.scala 96:25:@28503.4 package.scala 96:25:@28504.4]
  wire  x247; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 211:24:@28516.4]
  wire  _T_717; // @[FixedPoint.scala 50:25:@28523.4]
  wire [15:0] _T_721; // @[Bitwise.scala 72:12:@28525.4]
  wire [15:0] _T_722; // @[FixedPoint.scala 18:52:@28526.4]
  wire  _T_728; // @[Math.scala 451:55:@28528.4]
  wire [15:0] _T_729; // @[FixedPoint.scala 18:52:@28529.4]
  wire  _T_735; // @[Math.scala 451:110:@28531.4]
  wire  _T_736; // @[Math.scala 451:94:@28532.4]
  wire [31:0] _T_738; // @[Cat.scala 30:58:@28534.4]
  wire [31:0] _T_750; // @[Math.scala 406:56:@28544.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@28545.4]
  wire [31:0] x423_sum_number; // @[Math.scala 154:22:@28556.4 Math.scala 155:14:@28557.4]
  wire  _T_758; // @[FixedPoint.scala 50:25:@28561.4]
  wire [7:0] _T_762; // @[Bitwise.scala 72:12:@28563.4]
  wire [23:0] _T_763; // @[FixedPoint.scala 18:52:@28564.4]
  wire  _T_769; // @[Math.scala 451:55:@28566.4]
  wire [7:0] _T_770; // @[FixedPoint.scala 18:52:@28567.4]
  wire  _T_776; // @[Math.scala 451:110:@28569.4]
  wire  _T_777; // @[Math.scala 451:94:@28570.4]
  wire [31:0] _T_781; // @[package.scala 96:25:@28578.4 package.scala 96:25:@28579.4]
  wire [31:0] _T_791; // @[Math.scala 406:49:@28587.4]
  wire [31:0] _T_793; // @[Math.scala 406:56:@28589.4]
  wire [31:0] _T_794; // @[Math.scala 406:56:@28590.4]
  wire [31:0] _T_798; // @[package.scala 96:25:@28598.4]
  wire [31:0] x426_sum_number; // @[Math.scala 154:22:@28610.4 Math.scala 155:14:@28611.4]
  wire  _T_805; // @[FixedPoint.scala 50:25:@28615.4]
  wire [3:0] _T_809; // @[Bitwise.scala 72:12:@28617.4]
  wire [27:0] _T_810; // @[FixedPoint.scala 18:52:@28618.4]
  wire  _T_816; // @[Math.scala 451:55:@28620.4]
  wire [3:0] _T_817; // @[FixedPoint.scala 18:52:@28621.4]
  wire  _T_823; // @[Math.scala 451:110:@28623.4]
  wire  _T_824; // @[Math.scala 451:94:@28624.4]
  wire [31:0] _T_826; // @[Cat.scala 30:58:@28626.4]
  wire [31:0] _T_836; // @[Math.scala 406:49:@28634.4]
  wire [31:0] _T_838; // @[Math.scala 406:56:@28636.4]
  wire [31:0] _T_839; // @[Math.scala 406:56:@28637.4]
  wire [31:0] x429_sum_number; // @[Math.scala 154:22:@28648.4 Math.scala 155:14:@28649.4]
  wire  _T_846; // @[FixedPoint.scala 50:25:@28653.4]
  wire [1:0] _T_850; // @[Bitwise.scala 72:12:@28655.4]
  wire [29:0] _T_851; // @[FixedPoint.scala 18:52:@28656.4]
  wire  _T_857; // @[Math.scala 451:55:@28658.4]
  wire [1:0] _T_858; // @[FixedPoint.scala 18:52:@28659.4]
  wire  _T_864; // @[Math.scala 451:110:@28661.4]
  wire  _T_865; // @[Math.scala 451:94:@28662.4]
  wire [31:0] _T_867; // @[Cat.scala 30:58:@28664.4]
  wire [31:0] _T_877; // @[Math.scala 406:49:@28672.4]
  wire [31:0] _T_879; // @[Math.scala 406:56:@28674.4]
  wire [31:0] _T_880; // @[Math.scala 406:56:@28675.4]
  wire [31:0] x432_sum_number; // @[Math.scala 154:22:@28686.4 Math.scala 155:14:@28687.4]
  wire  _T_887; // @[FixedPoint.scala 50:25:@28691.4]
  wire [1:0] _T_891; // @[Bitwise.scala 72:12:@28693.4]
  wire [29:0] _T_892; // @[FixedPoint.scala 18:52:@28694.4]
  wire  _T_898; // @[Math.scala 451:55:@28696.4]
  wire [1:0] _T_899; // @[FixedPoint.scala 18:52:@28697.4]
  wire  _T_905; // @[Math.scala 451:110:@28699.4]
  wire  _T_906; // @[Math.scala 451:94:@28700.4]
  wire [31:0] _T_908; // @[Cat.scala 30:58:@28702.4]
  wire [31:0] _T_918; // @[Math.scala 406:49:@28710.4]
  wire [31:0] _T_920; // @[Math.scala 406:56:@28712.4]
  wire [31:0] _T_921; // @[Math.scala 406:56:@28713.4]
  wire [31:0] x435_sum_number; // @[Math.scala 154:22:@28724.4 Math.scala 155:14:@28725.4]
  wire  _T_928; // @[FixedPoint.scala 50:25:@28729.4]
  wire [1:0] _T_932; // @[Bitwise.scala 72:12:@28731.4]
  wire [29:0] _T_933; // @[FixedPoint.scala 18:52:@28732.4]
  wire  _T_939; // @[Math.scala 451:55:@28734.4]
  wire [1:0] _T_940; // @[FixedPoint.scala 18:52:@28735.4]
  wire  _T_946; // @[Math.scala 451:110:@28737.4]
  wire  _T_947; // @[Math.scala 451:94:@28738.4]
  wire [31:0] _T_949; // @[Cat.scala 30:58:@28740.4]
  wire [31:0] _T_959; // @[Math.scala 406:49:@28748.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@28750.4]
  wire [31:0] _T_962; // @[Math.scala 406:56:@28751.4]
  wire [31:0] x438_sum_number; // @[Math.scala 154:22:@28762.4 Math.scala 155:14:@28763.4]
  wire [31:0] _T_972; // @[Math.scala 476:37:@28768.4]
  wire  x439; // @[package.scala 96:25:@28776.4 package.scala 96:25:@28777.4]
  wire [31:0] x499_x438_sum_D1_number; // @[package.scala 96:25:@28811.4 package.scala 96:25:@28812.4]
  wire [31:0] x441_sub_number; // @[Math.scala 195:22:@28802.4 Math.scala 196:14:@28803.4]
  wire  _T_1029; // @[package.scala 96:25:@28875.4 package.scala 96:25:@28876.4]
  wire  _T_1031; // @[implicits.scala 55:10:@28877.4]
  wire  _T_1032; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 274:194:@28878.4]
  wire  x501_x248_D20; // @[package.scala 96:25:@28854.4 package.scala 96:25:@28855.4]
  wire  _T_1033; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 274:283:@28879.4]
  wire  _T_1034; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 274:291:@28880.4]
  wire [31:0] x254_rdcol_number; // @[Math.scala 195:22:@28899.4 Math.scala 196:14:@28900.4]
  wire [31:0] _T_1049; // @[Math.scala 476:37:@28905.4]
  wire  x255; // @[package.scala 96:25:@28913.4 package.scala 96:25:@28914.4]
  wire  x256; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 288:59:@28917.4]
  wire  _T_1062; // @[FixedPoint.scala 50:25:@28926.4]
  wire [15:0] _T_1066; // @[Bitwise.scala 72:12:@28928.4]
  wire [15:0] _T_1067; // @[FixedPoint.scala 18:52:@28929.4]
  wire  _T_1073; // @[Math.scala 451:55:@28931.4]
  wire [15:0] _T_1074; // @[FixedPoint.scala 18:52:@28932.4]
  wire  _T_1080; // @[Math.scala 451:110:@28934.4]
  wire  _T_1081; // @[Math.scala 451:94:@28935.4]
  wire [31:0] _T_1083; // @[Cat.scala 30:58:@28937.4]
  wire [31:0] _T_1095; // @[Math.scala 406:56:@28947.4]
  wire [31:0] _T_1096; // @[Math.scala 406:56:@28948.4]
  wire [31:0] x445_sum_number; // @[Math.scala 154:22:@28959.4 Math.scala 155:14:@28960.4]
  wire  _T_1103; // @[FixedPoint.scala 50:25:@28964.4]
  wire [7:0] _T_1107; // @[Bitwise.scala 72:12:@28966.4]
  wire [23:0] _T_1108; // @[FixedPoint.scala 18:52:@28967.4]
  wire  _T_1114; // @[Math.scala 451:55:@28969.4]
  wire [7:0] _T_1115; // @[FixedPoint.scala 18:52:@28970.4]
  wire  _T_1121; // @[Math.scala 451:110:@28972.4]
  wire  _T_1122; // @[Math.scala 451:94:@28973.4]
  wire [31:0] _T_1126; // @[package.scala 96:25:@28981.4 package.scala 96:25:@28982.4]
  wire [31:0] _T_1136; // @[Math.scala 406:49:@28990.4]
  wire [31:0] _T_1138; // @[Math.scala 406:56:@28992.4]
  wire [31:0] _T_1139; // @[Math.scala 406:56:@28993.4]
  wire [31:0] _T_1143; // @[package.scala 96:25:@29001.4]
  wire [31:0] x448_sum_number; // @[Math.scala 154:22:@29013.4 Math.scala 155:14:@29014.4]
  wire  _T_1150; // @[FixedPoint.scala 50:25:@29018.4]
  wire [3:0] _T_1154; // @[Bitwise.scala 72:12:@29020.4]
  wire [27:0] _T_1155; // @[FixedPoint.scala 18:52:@29021.4]
  wire  _T_1161; // @[Math.scala 451:55:@29023.4]
  wire [3:0] _T_1162; // @[FixedPoint.scala 18:52:@29024.4]
  wire  _T_1168; // @[Math.scala 451:110:@29026.4]
  wire  _T_1169; // @[Math.scala 451:94:@29027.4]
  wire [31:0] _T_1171; // @[Cat.scala 30:58:@29029.4]
  wire [31:0] _T_1181; // @[Math.scala 406:49:@29037.4]
  wire [31:0] _T_1183; // @[Math.scala 406:56:@29039.4]
  wire [31:0] _T_1184; // @[Math.scala 406:56:@29040.4]
  wire [31:0] x451_sum_number; // @[Math.scala 154:22:@29051.4 Math.scala 155:14:@29052.4]
  wire  _T_1191; // @[FixedPoint.scala 50:25:@29056.4]
  wire [1:0] _T_1195; // @[Bitwise.scala 72:12:@29058.4]
  wire [29:0] _T_1196; // @[FixedPoint.scala 18:52:@29059.4]
  wire  _T_1202; // @[Math.scala 451:55:@29061.4]
  wire [1:0] _T_1203; // @[FixedPoint.scala 18:52:@29062.4]
  wire  _T_1209; // @[Math.scala 451:110:@29064.4]
  wire  _T_1210; // @[Math.scala 451:94:@29065.4]
  wire [31:0] _T_1212; // @[Cat.scala 30:58:@29067.4]
  wire [31:0] _T_1222; // @[Math.scala 406:49:@29075.4]
  wire [31:0] _T_1224; // @[Math.scala 406:56:@29077.4]
  wire [31:0] _T_1225; // @[Math.scala 406:56:@29078.4]
  wire [31:0] x454_sum_number; // @[Math.scala 154:22:@29089.4 Math.scala 155:14:@29090.4]
  wire  _T_1232; // @[FixedPoint.scala 50:25:@29094.4]
  wire [1:0] _T_1236; // @[Bitwise.scala 72:12:@29096.4]
  wire [29:0] _T_1237; // @[FixedPoint.scala 18:52:@29097.4]
  wire  _T_1243; // @[Math.scala 451:55:@29099.4]
  wire [1:0] _T_1244; // @[FixedPoint.scala 18:52:@29100.4]
  wire  _T_1250; // @[Math.scala 451:110:@29102.4]
  wire  _T_1251; // @[Math.scala 451:94:@29103.4]
  wire [31:0] _T_1253; // @[Cat.scala 30:58:@29105.4]
  wire [31:0] _T_1263; // @[Math.scala 406:49:@29113.4]
  wire [31:0] _T_1265; // @[Math.scala 406:56:@29115.4]
  wire [31:0] _T_1266; // @[Math.scala 406:56:@29116.4]
  wire [31:0] x457_sum_number; // @[Math.scala 154:22:@29127.4 Math.scala 155:14:@29128.4]
  wire  _T_1273; // @[FixedPoint.scala 50:25:@29132.4]
  wire [1:0] _T_1277; // @[Bitwise.scala 72:12:@29134.4]
  wire [29:0] _T_1278; // @[FixedPoint.scala 18:52:@29135.4]
  wire  _T_1284; // @[Math.scala 451:55:@29137.4]
  wire [1:0] _T_1285; // @[FixedPoint.scala 18:52:@29138.4]
  wire  _T_1291; // @[Math.scala 451:110:@29140.4]
  wire  _T_1292; // @[Math.scala 451:94:@29141.4]
  wire [31:0] _T_1294; // @[Cat.scala 30:58:@29143.4]
  wire [31:0] _T_1304; // @[Math.scala 406:49:@29151.4]
  wire [31:0] _T_1306; // @[Math.scala 406:56:@29153.4]
  wire [31:0] _T_1307; // @[Math.scala 406:56:@29154.4]
  wire [31:0] x460_sum_number; // @[Math.scala 154:22:@29165.4 Math.scala 155:14:@29166.4]
  wire [31:0] _T_1317; // @[Math.scala 476:37:@29171.4]
  wire  x461; // @[package.scala 96:25:@29179.4 package.scala 96:25:@29180.4]
  wire [31:0] x503_x460_sum_D1_number; // @[package.scala 96:25:@29214.4 package.scala 96:25:@29215.4]
  wire [31:0] x463_sub_number; // @[Math.scala 195:22:@29205.4 Math.scala 196:14:@29206.4]
  wire  _T_1371; // @[package.scala 96:25:@29269.4 package.scala 96:25:@29270.4]
  wire  _T_1373; // @[implicits.scala 55:10:@29271.4]
  wire  _T_1374; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 351:194:@29272.4]
  wire  x504_x257_D20; // @[package.scala 96:25:@29248.4 package.scala 96:25:@29249.4]
  wire  _T_1375; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 351:283:@29273.4]
  wire  _T_1376; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 351:291:@29274.4]
  wire [31:0] x263_rdrow_number; // @[Math.scala 195:22:@29293.4 Math.scala 196:14:@29294.4]
  wire [31:0] _T_1393; // @[Math.scala 406:49:@29300.4]
  wire [31:0] _T_1395; // @[Math.scala 406:56:@29302.4]
  wire [31:0] _T_1396; // @[Math.scala 406:56:@29303.4]
  wire [31:0] x465_number; // @[implicits.scala 133:21:@29304.4]
  wire  x265; // @[package.scala 96:25:@29318.4 package.scala 96:25:@29319.4]
  wire  x506_x240_D1; // @[package.scala 96:25:@29327.4 package.scala 96:25:@29328.4]
  wire  x266; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 363:24:@29331.4]
  wire [31:0] _T_1422; // @[Math.scala 406:49:@29340.4]
  wire [31:0] _T_1424; // @[Math.scala 406:56:@29342.4]
  wire [31:0] _T_1425; // @[Math.scala 406:56:@29343.4]
  wire [31:0] _T_1429; // @[package.scala 96:25:@29351.4]
  wire  _T_1433; // @[FixedPoint.scala 50:25:@29358.4]
  wire [1:0] _T_1437; // @[Bitwise.scala 72:12:@29360.4]
  wire [29:0] _T_1438; // @[FixedPoint.scala 18:52:@29361.4]
  wire  _T_1444; // @[Math.scala 451:55:@29363.4]
  wire [1:0] _T_1445; // @[FixedPoint.scala 18:52:@29364.4]
  wire  _T_1451; // @[Math.scala 451:110:@29366.4]
  wire  _T_1452; // @[Math.scala 451:94:@29367.4]
  wire [31:0] _T_1456; // @[package.scala 96:25:@29375.4 package.scala 96:25:@29376.4]
  wire [31:0] x269_1_number; // @[Math.scala 454:20:@29377.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@29382.4]
  wire [40:0] _T_1461; // @[Math.scala 461:32:@29382.4]
  wire [38:0] _GEN_3; // @[Math.scala 461:32:@29387.4]
  wire [38:0] _T_1464; // @[Math.scala 461:32:@29387.4]
  wire  _T_1497; // @[package.scala 96:25:@29464.4 package.scala 96:25:@29465.4]
  wire  _T_1499; // @[implicits.scala 55:10:@29466.4]
  wire  _T_1500; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 392:194:@29467.4]
  wire  x511_x267_D20; // @[package.scala 96:25:@29452.4 package.scala 96:25:@29453.4]
  wire  _T_1501; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 392:283:@29468.4]
  wire  _T_1502; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 392:291:@29469.4]
  wire  x274; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 402:59:@29480.4]
  wire  _T_1531; // @[package.scala 96:25:@29524.4 package.scala 96:25:@29525.4]
  wire  _T_1533; // @[implicits.scala 55:10:@29526.4]
  wire  _T_1534; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 417:194:@29527.4]
  wire  x513_x275_D20; // @[package.scala 96:25:@29512.4 package.scala 96:25:@29513.4]
  wire  _T_1535; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 417:283:@29528.4]
  wire  _T_1536; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 417:291:@29529.4]
  wire  x279; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 421:59:@29540.4]
  wire  _T_1560; // @[package.scala 96:25:@29573.4 package.scala 96:25:@29574.4]
  wire  _T_1562; // @[implicits.scala 55:10:@29575.4]
  wire  _T_1563; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 432:194:@29576.4]
  wire  x514_x280_D20; // @[package.scala 96:25:@29561.4 package.scala 96:25:@29562.4]
  wire  _T_1564; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 432:283:@29577.4]
  wire  _T_1565; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 432:291:@29578.4]
  wire [31:0] x284_rdrow_number; // @[Math.scala 195:22:@29597.4 Math.scala 196:14:@29598.4]
  wire [31:0] _T_1582; // @[Math.scala 406:49:@29604.4]
  wire [31:0] _T_1584; // @[Math.scala 406:56:@29606.4]
  wire [31:0] _T_1585; // @[Math.scala 406:56:@29607.4]
  wire [31:0] x470_number; // @[implicits.scala 133:21:@29608.4]
  wire  x286; // @[package.scala 96:25:@29622.4 package.scala 96:25:@29623.4]
  wire  x287; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 442:24:@29626.4]
  wire [31:0] _T_1608; // @[Math.scala 406:49:@29635.4]
  wire [31:0] _T_1610; // @[Math.scala 406:56:@29637.4]
  wire [31:0] _T_1611; // @[Math.scala 406:56:@29638.4]
  wire [31:0] _T_1615; // @[package.scala 96:25:@29646.4]
  wire  _T_1619; // @[FixedPoint.scala 50:25:@29653.4]
  wire [1:0] _T_1623; // @[Bitwise.scala 72:12:@29655.4]
  wire [29:0] _T_1624; // @[FixedPoint.scala 18:52:@29656.4]
  wire  _T_1630; // @[Math.scala 451:55:@29658.4]
  wire [1:0] _T_1631; // @[FixedPoint.scala 18:52:@29659.4]
  wire  _T_1637; // @[Math.scala 451:110:@29661.4]
  wire  _T_1638; // @[Math.scala 451:94:@29662.4]
  wire [31:0] _T_1642; // @[package.scala 96:25:@29670.4 package.scala 96:25:@29671.4]
  wire [31:0] x290_1_number; // @[Math.scala 454:20:@29672.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@29677.4]
  wire [40:0] _T_1647; // @[Math.scala 461:32:@29677.4]
  wire [38:0] _GEN_5; // @[Math.scala 461:32:@29682.4]
  wire [38:0] _T_1650; // @[Math.scala 461:32:@29682.4]
  wire  _T_1680; // @[package.scala 96:25:@29750.4 package.scala 96:25:@29751.4]
  wire  _T_1682; // @[implicits.scala 55:10:@29752.4]
  wire  _T_1683; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 469:194:@29753.4]
  wire  x516_x288_D20; // @[package.scala 96:25:@29720.4 package.scala 96:25:@29721.4]
  wire  _T_1684; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 469:283:@29754.4]
  wire  _T_1685; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 469:291:@29755.4]
  wire  x295; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 473:24:@29766.4]
  wire  _T_1712; // @[package.scala 96:25:@29808.4 package.scala 96:25:@29809.4]
  wire  _T_1714; // @[implicits.scala 55:10:@29810.4]
  wire  _T_1715; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 486:194:@29811.4]
  wire  x520_x296_D20; // @[package.scala 96:25:@29796.4 package.scala 96:25:@29797.4]
  wire  _T_1716; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 486:283:@29812.4]
  wire  _T_1717; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 486:291:@29813.4]
  wire  x300; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 490:24:@29824.4]
  wire  _T_1741; // @[package.scala 96:25:@29857.4 package.scala 96:25:@29858.4]
  wire  _T_1743; // @[implicits.scala 55:10:@29859.4]
  wire  _T_1744; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 501:194:@29860.4]
  wire  x521_x301_D20; // @[package.scala 96:25:@29845.4 package.scala 96:25:@29846.4]
  wire  _T_1745; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 501:283:@29861.4]
  wire  _T_1746; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 501:291:@29862.4]
  wire [31:0] x325_sub_number; // @[Math.scala 195:22:@30117.4 Math.scala 196:14:@30118.4]
  wire [31:0] x327_sub_number; // @[Math.scala 195:22:@30139.4 Math.scala 196:14:@30140.4]
  wire  x326; // @[package.scala 96:25:@30129.4 package.scala 96:25:@30130.4]
  wire  x328; // @[package.scala 96:25:@30151.4 package.scala 96:25:@30152.4]
  wire  x329; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 565:24:@30155.4]
  wire [31:0] x524_x325_sub_D1_number; // @[package.scala 96:25:@30163.4 package.scala 96:25:@30164.4]
  wire  _T_1928; // @[package.scala 96:25:@30257.4 package.scala 96:25:@30258.4]
  wire  _T_1930; // @[implicits.scala 55:10:@30259.4]
  wire  x526_b223_D75; // @[package.scala 96:25:@30239.4 package.scala 96:25:@30240.4]
  wire  _T_1931; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 589:117:@30260.4]
  wire  x527_b224_D75; // @[package.scala 96:25:@30248.4 package.scala 96:25:@30249.4]
  wire  _T_1932; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 589:123:@30261.4]
  wire [31:0] x236_sum_number; // @[Math.scala 154:22:@28277.4 Math.scala 155:14:@28278.4]
  wire [31:0] x485_x417_D13_number; // @[package.scala 96:25:@28286.4 package.scala 96:25:@28287.4]
  wire [31:0] x489_x395_D21_number; // @[package.scala 96:25:@28322.4 package.scala 96:25:@28323.4]
  wire [31:0] x492_x417_D37_number; // @[package.scala 96:25:@28408.4 package.scala 96:25:@28409.4]
  wire [31:0] x494_x236_sum_D24_number; // @[package.scala 96:25:@28426.4 package.scala 96:25:@28427.4]
  wire [31:0] x497_x395_D45_number; // @[package.scala 96:25:@28453.4 package.scala 96:25:@28454.4]
  wire [31:0] x251_sum_number; // @[Math.scala 154:22:@28845.4 Math.scala 155:14:@28846.4]
  wire [31:0] x502_x442_D13_number; // @[package.scala 96:25:@28863.4 package.scala 96:25:@28864.4]
  wire [31:0] x260_sum_number; // @[Math.scala 154:22:@29239.4 Math.scala 155:14:@29240.4]
  wire [31:0] x505_x464_D13_number; // @[package.scala 96:25:@29257.4 package.scala 96:25:@29258.4]
  wire [31:0] x509_x466_D20_number; // @[package.scala 96:25:@29434.4 package.scala 96:25:@29435.4]
  wire [31:0] x510_x271_sum_D1_number; // @[package.scala 96:25:@29443.4 package.scala 96:25:@29444.4]
  wire [31:0] x276_sum_number; // @[Math.scala 154:22:@29503.4 Math.scala 155:14:@29504.4]
  wire [31:0] x281_sum_number; // @[Math.scala 154:22:@29552.4 Math.scala 155:14:@29553.4]
  wire [31:0] x517_x292_sum_D1_number; // @[package.scala 96:25:@29729.4 package.scala 96:25:@29730.4]
  wire [31:0] x518_x471_D20_number; // @[package.scala 96:25:@29738.4 package.scala 96:25:@29739.4]
  wire [31:0] x297_sum_number; // @[Math.scala 154:22:@29787.4 Math.scala 155:14:@29788.4]
  wire [31:0] x302_sum_number; // @[Math.scala 154:22:@29836.4 Math.scala 155:14:@29837.4]
  _ _ ( // @[Math.scala 720:24:@27771.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@27783.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@27806.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x227_lb_0 x227_lb_0 ( // @[m_x227_lb_0.scala 35:17:@27816.4]
    .clock(x227_lb_0_clock),
    .reset(x227_lb_0_reset),
    .io_rPort_8_banks_1(x227_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x227_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x227_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x227_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x227_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x227_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x227_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x227_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x227_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x227_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x227_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x227_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x227_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x227_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x227_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x227_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x227_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x227_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x227_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x227_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x227_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x227_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x227_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x227_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x227_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x227_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x227_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x227_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x227_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x227_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x227_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x227_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x227_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x227_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x227_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x227_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x227_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x227_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x227_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x227_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x227_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x227_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x227_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x227_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x227_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x227_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x227_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x227_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x227_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x227_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x227_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x227_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x227_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x227_lb_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x227_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x227_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x227_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x227_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x227_lb_0_io_wPort_0_en_0)
  );
  x208_sum x398_sum_1 ( // @[Math.scala 150:24:@27941.4]
    .clock(x398_sum_1_clock),
    .reset(x398_sum_1_reset),
    .io_a(x398_sum_1_io_a),
    .io_b(x398_sum_1_io_b),
    .io_flow(x398_sum_1_io_flow),
    .io_result(x398_sum_1_io_result)
  );
  x208_sum x401_sum_1 ( // @[Math.scala 150:24:@27979.4]
    .clock(x401_sum_1_clock),
    .reset(x401_sum_1_reset),
    .io_a(x401_sum_1_io_a),
    .io_b(x401_sum_1_io_b),
    .io_flow(x401_sum_1_io_flow),
    .io_result(x401_sum_1_io_result)
  );
  x208_sum x404_sum_1 ( // @[Math.scala 150:24:@28017.4]
    .clock(x404_sum_1_clock),
    .reset(x404_sum_1_reset),
    .io_a(x404_sum_1_io_a),
    .io_b(x404_sum_1_io_b),
    .io_flow(x404_sum_1_io_flow),
    .io_result(x404_sum_1_io_result)
  );
  x208_sum x407_sum_1 ( // @[Math.scala 150:24:@28055.4]
    .clock(x407_sum_1_clock),
    .reset(x407_sum_1_reset),
    .io_a(x407_sum_1_io_a),
    .io_b(x407_sum_1_io_b),
    .io_flow(x407_sum_1_io_flow),
    .io_result(x407_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@28078.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_2 ( // @[package.scala 93:22:@28096.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x208_sum x410_sum_1 ( // @[Math.scala 150:24:@28109.4]
    .clock(x410_sum_1_clock),
    .reset(x410_sum_1_reset),
    .io_a(x410_sum_1_io_a),
    .io_b(x410_sum_1_io_b),
    .io_flow(x410_sum_1_io_flow),
    .io_result(x410_sum_1_io_result)
  );
  x208_sum x413_sum_1 ( // @[Math.scala 150:24:@28147.4]
    .clock(x413_sum_1_clock),
    .reset(x413_sum_1_reset),
    .io_a(x413_sum_1_io_a),
    .io_b(x413_sum_1_io_b),
    .io_flow(x413_sum_1_io_flow),
    .io_result(x413_sum_1_io_result)
  );
  x390_sub x416_sub_1 ( // @[Math.scala 191:24:@28173.4]
    .clock(x416_sub_1_clock),
    .reset(x416_sub_1_reset),
    .io_a(x416_sub_1_io_a),
    .io_b(x416_sub_1_io_b),
    .io_flow(x416_sub_1_io_flow),
    .io_result(x416_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@28183.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@28192.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_5 ( // @[package.scala 93:22:@28201.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x208_sum x420_sum_1 ( // @[Math.scala 150:24:@28240.4]
    .clock(x420_sum_1_clock),
    .reset(x420_sum_1_reset),
    .io_a(x420_sum_1_io_a),
    .io_b(x420_sum_1_io_b),
    .io_flow(x420_sum_1_io_flow),
    .io_result(x420_sum_1_io_result)
  );
  x235_div x235_div_1 ( // @[Math.scala 327:24:@28252.4]
    .clock(x235_div_1_clock),
    .io_a(x235_div_1_io_a),
    .io_flow(x235_div_1_io_flow),
    .io_result(x235_div_1_io_result)
  );
  RetimeWrapper_184 RetimeWrapper_6 ( // @[package.scala 93:22:@28262.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x208_sum x236_sum_1 ( // @[Math.scala 150:24:@28271.4]
    .clock(x236_sum_1_clock),
    .reset(x236_sum_1_reset),
    .io_a(x236_sum_1_io_a),
    .io_b(x236_sum_1_io_b),
    .io_flow(x236_sum_1_io_flow),
    .io_result(x236_sum_1_io_result)
  );
  RetimeWrapper_186 RetimeWrapper_7 ( // @[package.scala 93:22:@28281.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_8 ( // @[package.scala 93:22:@28290.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_9 ( // @[package.scala 93:22:@28299.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_10 ( // @[package.scala 93:22:@28308.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_190 RetimeWrapper_11 ( // @[package.scala 93:22:@28317.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_12 ( // @[package.scala 93:22:@28328.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_192 RetimeWrapper_13 ( // @[package.scala 93:22:@28349.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@28363.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_192 RetimeWrapper_15 ( // @[package.scala 93:22:@28372.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@28388.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_196 RetimeWrapper_17 ( // @[package.scala 93:22:@28403.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_18 ( // @[package.scala 93:22:@28412.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_19 ( // @[package.scala 93:22:@28421.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_20 ( // @[package.scala 93:22:@28430.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_21 ( // @[package.scala 93:22:@28439.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_22 ( // @[package.scala 93:22:@28448.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_23 ( // @[package.scala 93:22:@28460.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  x390_sub x245_rdcol_1 ( // @[Math.scala 191:24:@28483.4]
    .clock(x245_rdcol_1_clock),
    .reset(x245_rdcol_1_reset),
    .io_a(x245_rdcol_1_io_a),
    .io_b(x245_rdcol_1_io_b),
    .io_flow(x245_rdcol_1_io_flow),
    .io_result(x245_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@28498.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@28507.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  x208_sum x423_sum_1 ( // @[Math.scala 150:24:@28550.4]
    .clock(x423_sum_1_clock),
    .reset(x423_sum_1_reset),
    .io_a(x423_sum_1_io_a),
    .io_b(x423_sum_1_io_b),
    .io_flow(x423_sum_1_io_flow),
    .io_result(x423_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_26 ( // @[package.scala 93:22:@28573.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_27 ( // @[package.scala 93:22:@28591.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x208_sum x426_sum_1 ( // @[Math.scala 150:24:@28604.4]
    .clock(x426_sum_1_clock),
    .reset(x426_sum_1_reset),
    .io_a(x426_sum_1_io_a),
    .io_b(x426_sum_1_io_b),
    .io_flow(x426_sum_1_io_flow),
    .io_result(x426_sum_1_io_result)
  );
  x208_sum x429_sum_1 ( // @[Math.scala 150:24:@28642.4]
    .clock(x429_sum_1_clock),
    .reset(x429_sum_1_reset),
    .io_a(x429_sum_1_io_a),
    .io_b(x429_sum_1_io_b),
    .io_flow(x429_sum_1_io_flow),
    .io_result(x429_sum_1_io_result)
  );
  x208_sum x432_sum_1 ( // @[Math.scala 150:24:@28680.4]
    .clock(x432_sum_1_clock),
    .reset(x432_sum_1_reset),
    .io_a(x432_sum_1_io_a),
    .io_b(x432_sum_1_io_b),
    .io_flow(x432_sum_1_io_flow),
    .io_result(x432_sum_1_io_result)
  );
  x208_sum x435_sum_1 ( // @[Math.scala 150:24:@28718.4]
    .clock(x435_sum_1_clock),
    .reset(x435_sum_1_reset),
    .io_a(x435_sum_1_io_a),
    .io_b(x435_sum_1_io_b),
    .io_flow(x435_sum_1_io_flow),
    .io_result(x435_sum_1_io_result)
  );
  x208_sum x438_sum_1 ( // @[Math.scala 150:24:@28756.4]
    .clock(x438_sum_1_clock),
    .reset(x438_sum_1_reset),
    .io_a(x438_sum_1_io_a),
    .io_b(x438_sum_1_io_b),
    .io_flow(x438_sum_1_io_flow),
    .io_result(x438_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@28771.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@28785.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  x390_sub x441_sub_1 ( // @[Math.scala 191:24:@28796.4]
    .clock(x441_sub_1_clock),
    .reset(x441_sub_1_reset),
    .io_a(x441_sub_1_io_a),
    .io_b(x441_sub_1_io_b),
    .io_flow(x441_sub_1_io_flow),
    .io_result(x441_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_30 ( // @[package.scala 93:22:@28806.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x235_div x250_div_1 ( // @[Math.scala 327:24:@28820.4]
    .clock(x250_div_1_clock),
    .io_a(x250_div_1_io_a),
    .io_flow(x250_div_1_io_flow),
    .io_result(x250_div_1_io_result)
  );
  RetimeWrapper_218 RetimeWrapper_31 ( // @[package.scala 93:22:@28830.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x208_sum x251_sum_1 ( // @[Math.scala 150:24:@28839.4]
    .clock(x251_sum_1_clock),
    .reset(x251_sum_1_reset),
    .io_a(x251_sum_1_io_a),
    .io_b(x251_sum_1_io_b),
    .io_flow(x251_sum_1_io_flow),
    .io_result(x251_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_32 ( // @[package.scala 93:22:@28849.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_33 ( // @[package.scala 93:22:@28858.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_34 ( // @[package.scala 93:22:@28870.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x390_sub x254_rdcol_1 ( // @[Math.scala 191:24:@28893.4]
    .clock(x254_rdcol_1_clock),
    .reset(x254_rdcol_1_reset),
    .io_a(x254_rdcol_1_io_a),
    .io_b(x254_rdcol_1_io_b),
    .io_flow(x254_rdcol_1_io_flow),
    .io_result(x254_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@28908.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  x208_sum x445_sum_1 ( // @[Math.scala 150:24:@28953.4]
    .clock(x445_sum_1_clock),
    .reset(x445_sum_1_reset),
    .io_a(x445_sum_1_io_a),
    .io_b(x445_sum_1_io_b),
    .io_flow(x445_sum_1_io_flow),
    .io_result(x445_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_36 ( // @[package.scala 93:22:@28976.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_37 ( // @[package.scala 93:22:@28994.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x208_sum x448_sum_1 ( // @[Math.scala 150:24:@29007.4]
    .clock(x448_sum_1_clock),
    .reset(x448_sum_1_reset),
    .io_a(x448_sum_1_io_a),
    .io_b(x448_sum_1_io_b),
    .io_flow(x448_sum_1_io_flow),
    .io_result(x448_sum_1_io_result)
  );
  x208_sum x451_sum_1 ( // @[Math.scala 150:24:@29045.4]
    .clock(x451_sum_1_clock),
    .reset(x451_sum_1_reset),
    .io_a(x451_sum_1_io_a),
    .io_b(x451_sum_1_io_b),
    .io_flow(x451_sum_1_io_flow),
    .io_result(x451_sum_1_io_result)
  );
  x208_sum x454_sum_1 ( // @[Math.scala 150:24:@29083.4]
    .clock(x454_sum_1_clock),
    .reset(x454_sum_1_reset),
    .io_a(x454_sum_1_io_a),
    .io_b(x454_sum_1_io_b),
    .io_flow(x454_sum_1_io_flow),
    .io_result(x454_sum_1_io_result)
  );
  x208_sum x457_sum_1 ( // @[Math.scala 150:24:@29121.4]
    .clock(x457_sum_1_clock),
    .reset(x457_sum_1_reset),
    .io_a(x457_sum_1_io_a),
    .io_b(x457_sum_1_io_b),
    .io_flow(x457_sum_1_io_flow),
    .io_result(x457_sum_1_io_result)
  );
  x208_sum x460_sum_1 ( // @[Math.scala 150:24:@29159.4]
    .clock(x460_sum_1_clock),
    .reset(x460_sum_1_reset),
    .io_a(x460_sum_1_io_a),
    .io_b(x460_sum_1_io_b),
    .io_flow(x460_sum_1_io_flow),
    .io_result(x460_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@29174.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper RetimeWrapper_39 ( // @[package.scala 93:22:@29188.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x390_sub x463_sub_1 ( // @[Math.scala 191:24:@29199.4]
    .clock(x463_sub_1_clock),
    .reset(x463_sub_1_reset),
    .io_a(x463_sub_1_io_a),
    .io_b(x463_sub_1_io_b),
    .io_flow(x463_sub_1_io_flow),
    .io_result(x463_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_40 ( // @[package.scala 93:22:@29209.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x235_div x259_div_1 ( // @[Math.scala 327:24:@29223.4]
    .clock(x259_div_1_clock),
    .io_a(x259_div_1_io_a),
    .io_flow(x259_div_1_io_flow),
    .io_result(x259_div_1_io_result)
  );
  x208_sum x260_sum_1 ( // @[Math.scala 150:24:@29233.4]
    .clock(x260_sum_1_clock),
    .reset(x260_sum_1_reset),
    .io_a(x260_sum_1_io_a),
    .io_b(x260_sum_1_io_b),
    .io_flow(x260_sum_1_io_flow),
    .io_result(x260_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_41 ( // @[package.scala 93:22:@29243.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_42 ( // @[package.scala 93:22:@29252.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_43 ( // @[package.scala 93:22:@29264.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x390_sub x263_rdrow_1 ( // @[Math.scala 191:24:@29287.4]
    .clock(x263_rdrow_1_clock),
    .reset(x263_rdrow_1_reset),
    .io_a(x263_rdrow_1_io_a),
    .io_b(x263_rdrow_1_io_b),
    .io_flow(x263_rdrow_1_io_flow),
    .io_result(x263_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@29313.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@29322.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_46 ( // @[package.scala 93:22:@29344.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_47 ( // @[package.scala 93:22:@29370.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  x208_sum x469_sum_1 ( // @[Math.scala 150:24:@29391.4]
    .clock(x469_sum_1_clock),
    .reset(x469_sum_1_reset),
    .io_a(x469_sum_1_io_a),
    .io_b(x469_sum_1_io_b),
    .io_flow(x469_sum_1_io_flow),
    .io_result(x469_sum_1_io_result)
  );
  RetimeWrapper_247 RetimeWrapper_48 ( // @[package.scala 93:22:@29401.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_192 RetimeWrapper_49 ( // @[package.scala 93:22:@29410.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  x208_sum x271_sum_1 ( // @[Math.scala 150:24:@29419.4]
    .clock(x271_sum_1_clock),
    .reset(x271_sum_1_reset),
    .io_a(x271_sum_1_io_a),
    .io_b(x271_sum_1_io_b),
    .io_flow(x271_sum_1_io_flow),
    .io_result(x271_sum_1_io_result)
  );
  RetimeWrapper_188 RetimeWrapper_50 ( // @[package.scala 93:22:@29429.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_51 ( // @[package.scala 93:22:@29438.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_52 ( // @[package.scala 93:22:@29447.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_53 ( // @[package.scala 93:22:@29459.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_254 RetimeWrapper_54 ( // @[package.scala 93:22:@29486.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x208_sum x276_sum_1 ( // @[Math.scala 150:24:@29497.4]
    .clock(x276_sum_1_clock),
    .reset(x276_sum_1_reset),
    .io_a(x276_sum_1_io_a),
    .io_b(x276_sum_1_io_b),
    .io_flow(x276_sum_1_io_flow),
    .io_result(x276_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_55 ( // @[package.scala 93:22:@29507.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_56 ( // @[package.scala 93:22:@29519.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x208_sum x281_sum_1 ( // @[Math.scala 150:24:@29546.4]
    .clock(x281_sum_1_clock),
    .reset(x281_sum_1_reset),
    .io_a(x281_sum_1_io_a),
    .io_b(x281_sum_1_io_b),
    .io_flow(x281_sum_1_io_flow),
    .io_result(x281_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_57 ( // @[package.scala 93:22:@29556.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_58 ( // @[package.scala 93:22:@29568.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x390_sub x284_rdrow_1 ( // @[Math.scala 191:24:@29591.4]
    .clock(x284_rdrow_1_clock),
    .reset(x284_rdrow_1_reset),
    .io_a(x284_rdrow_1_io_a),
    .io_b(x284_rdrow_1_io_b),
    .io_flow(x284_rdrow_1_io_flow),
    .io_result(x284_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_59 ( // @[package.scala 93:22:@29617.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_60 ( // @[package.scala 93:22:@29639.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_61 ( // @[package.scala 93:22:@29665.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x208_sum x474_sum_1 ( // @[Math.scala 150:24:@29686.4]
    .clock(x474_sum_1_clock),
    .reset(x474_sum_1_reset),
    .io_a(x474_sum_1_io_a),
    .io_b(x474_sum_1_io_b),
    .io_flow(x474_sum_1_io_flow),
    .io_result(x474_sum_1_io_result)
  );
  RetimeWrapper_247 RetimeWrapper_62 ( // @[package.scala 93:22:@29696.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x208_sum x292_sum_1 ( // @[Math.scala 150:24:@29705.4]
    .clock(x292_sum_1_clock),
    .reset(x292_sum_1_reset),
    .io_a(x292_sum_1_io_a),
    .io_b(x292_sum_1_io_b),
    .io_flow(x292_sum_1_io_flow),
    .io_result(x292_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_63 ( // @[package.scala 93:22:@29715.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_64 ( // @[package.scala 93:22:@29724.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_65 ( // @[package.scala 93:22:@29733.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_66 ( // @[package.scala 93:22:@29745.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_254 RetimeWrapper_67 ( // @[package.scala 93:22:@29772.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x208_sum x297_sum_1 ( // @[Math.scala 150:24:@29781.4]
    .clock(x297_sum_1_clock),
    .reset(x297_sum_1_reset),
    .io_a(x297_sum_1_io_a),
    .io_b(x297_sum_1_io_b),
    .io_flow(x297_sum_1_io_flow),
    .io_result(x297_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_68 ( // @[package.scala 93:22:@29791.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_69 ( // @[package.scala 93:22:@29803.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x208_sum x302_sum_1 ( // @[Math.scala 150:24:@29830.4]
    .clock(x302_sum_1_clock),
    .reset(x302_sum_1_reset),
    .io_a(x302_sum_1_io_a),
    .io_b(x302_sum_1_io_b),
    .io_flow(x302_sum_1_io_flow),
    .io_result(x302_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_70 ( // @[package.scala 93:22:@29840.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_71 ( // @[package.scala 93:22:@29852.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x305 x305_1 ( // @[Math.scala 262:24:@29875.4]
    .clock(x305_1_clock),
    .io_a(x305_1_io_a),
    .io_b(x305_1_io_b),
    .io_flow(x305_1_io_flow),
    .io_result(x305_1_io_result)
  );
  x305 x306_1 ( // @[Math.scala 262:24:@29887.4]
    .clock(x306_1_clock),
    .io_a(x306_1_io_a),
    .io_b(x306_1_io_b),
    .io_flow(x306_1_io_flow),
    .io_result(x306_1_io_result)
  );
  x305 x307_1 ( // @[Math.scala 262:24:@29899.4]
    .clock(x307_1_clock),
    .io_a(x307_1_io_a),
    .io_b(x307_1_io_b),
    .io_flow(x307_1_io_flow),
    .io_result(x307_1_io_result)
  );
  x305 x308_1 ( // @[Math.scala 262:24:@29911.4]
    .clock(x308_1_clock),
    .io_a(x308_1_io_a),
    .io_b(x308_1_io_b),
    .io_flow(x308_1_io_flow),
    .io_result(x308_1_io_result)
  );
  x305 x309_1 ( // @[Math.scala 262:24:@29923.4]
    .clock(x309_1_clock),
    .io_a(x309_1_io_a),
    .io_b(x309_1_io_b),
    .io_flow(x309_1_io_flow),
    .io_result(x309_1_io_result)
  );
  x305 x310_1 ( // @[Math.scala 262:24:@29937.4]
    .clock(x310_1_clock),
    .io_a(x310_1_io_a),
    .io_b(x310_1_io_b),
    .io_flow(x310_1_io_flow),
    .io_result(x310_1_io_result)
  );
  x305 x311_1 ( // @[Math.scala 262:24:@29949.4]
    .clock(x311_1_clock),
    .io_a(x311_1_io_a),
    .io_b(x311_1_io_b),
    .io_flow(x311_1_io_flow),
    .io_result(x311_1_io_result)
  );
  x305 x312_1 ( // @[Math.scala 262:24:@29961.4]
    .clock(x312_1_clock),
    .io_a(x312_1_io_a),
    .io_b(x312_1_io_b),
    .io_flow(x312_1_io_flow),
    .io_result(x312_1_io_result)
  );
  x305 x313_1 ( // @[Math.scala 262:24:@29973.4]
    .clock(x313_1_clock),
    .io_a(x313_1_io_a),
    .io_b(x313_1_io_b),
    .io_flow(x313_1_io_flow),
    .io_result(x313_1_io_result)
  );
  x314_x13 x314_x13_1 ( // @[Math.scala 150:24:@29983.4]
    .clock(x314_x13_1_clock),
    .reset(x314_x13_1_reset),
    .io_a(x314_x13_1_io_a),
    .io_b(x314_x13_1_io_b),
    .io_flow(x314_x13_1_io_flow),
    .io_result(x314_x13_1_io_result)
  );
  x314_x13 x315_x14_1 ( // @[Math.scala 150:24:@29993.4]
    .clock(x315_x14_1_clock),
    .reset(x315_x14_1_reset),
    .io_a(x315_x14_1_io_a),
    .io_b(x315_x14_1_io_b),
    .io_flow(x315_x14_1_io_flow),
    .io_result(x315_x14_1_io_result)
  );
  x314_x13 x316_x13_1 ( // @[Math.scala 150:24:@30003.4]
    .clock(x316_x13_1_clock),
    .reset(x316_x13_1_reset),
    .io_a(x316_x13_1_io_a),
    .io_b(x316_x13_1_io_b),
    .io_flow(x316_x13_1_io_flow),
    .io_result(x316_x13_1_io_result)
  );
  x314_x13 x317_x14_1 ( // @[Math.scala 150:24:@30013.4]
    .clock(x317_x14_1_clock),
    .reset(x317_x14_1_reset),
    .io_a(x317_x14_1_io_a),
    .io_b(x317_x14_1_io_b),
    .io_flow(x317_x14_1_io_flow),
    .io_result(x317_x14_1_io_result)
  );
  x314_x13 x318_x13_1 ( // @[Math.scala 150:24:@30023.4]
    .clock(x318_x13_1_clock),
    .reset(x318_x13_1_reset),
    .io_a(x318_x13_1_io_a),
    .io_b(x318_x13_1_io_b),
    .io_flow(x318_x13_1_io_flow),
    .io_result(x318_x13_1_io_result)
  );
  x314_x13 x319_x14_1 ( // @[Math.scala 150:24:@30033.4]
    .clock(x319_x14_1_clock),
    .reset(x319_x14_1_reset),
    .io_a(x319_x14_1_io_a),
    .io_b(x319_x14_1_io_b),
    .io_flow(x319_x14_1_io_flow),
    .io_result(x319_x14_1_io_result)
  );
  x314_x13 x320_x13_1 ( // @[Math.scala 150:24:@30043.4]
    .clock(x320_x13_1_clock),
    .reset(x320_x13_1_reset),
    .io_a(x320_x13_1_io_a),
    .io_b(x320_x13_1_io_b),
    .io_flow(x320_x13_1_io_flow),
    .io_result(x320_x13_1_io_result)
  );
  RetimeWrapper_286 RetimeWrapper_72 ( // @[package.scala 93:22:@30053.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x314_x13 x321_sum_1 ( // @[Math.scala 150:24:@30062.4]
    .clock(x321_sum_1_clock),
    .reset(x321_sum_1_reset),
    .io_a(x321_sum_1_io_a),
    .io_b(x321_sum_1_io_b),
    .io_flow(x321_sum_1_io_flow),
    .io_result(x321_sum_1_io_result)
  );
  x322 x322_1 ( // @[Math.scala 720:24:@30072.4]
    .io_b(x322_1_io_b),
    .io_result(x322_1_io_result)
  );
  x323_mul x323_mul_1 ( // @[Math.scala 262:24:@30083.4]
    .clock(x323_mul_1_clock),
    .io_a(x323_mul_1_io_a),
    .io_b(x323_mul_1_io_b),
    .io_flow(x323_mul_1_io_flow),
    .io_result(x323_mul_1_io_result)
  );
  x324 x324_1 ( // @[Math.scala 720:24:@30093.4]
    .io_b(x324_1_io_b),
    .io_result(x324_1_io_result)
  );
  RetimeWrapper_288 RetimeWrapper_73 ( // @[package.scala 93:22:@30102.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x325_sub x325_sub_1 ( // @[Math.scala 191:24:@30111.4]
    .clock(x325_sub_1_clock),
    .reset(x325_sub_1_reset),
    .io_a(x325_sub_1_io_a),
    .io_b(x325_sub_1_io_b),
    .io_flow(x325_sub_1_io_flow),
    .io_result(x325_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_74 ( // @[package.scala 93:22:@30124.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x325_sub x327_sub_1 ( // @[Math.scala 191:24:@30133.4]
    .clock(x327_sub_1_clock),
    .reset(x327_sub_1_reset),
    .io_a(x327_sub_1_io_a),
    .io_b(x327_sub_1_io_b),
    .io_flow(x327_sub_1_io_flow),
    .io_result(x327_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_75 ( // @[package.scala 93:22:@30146.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_76 ( // @[package.scala 93:22:@30158.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x322 x331_1 ( // @[Math.scala 720:24:@30172.4]
    .io_b(x331_1_io_b),
    .io_result(x331_1_io_result)
  );
  x323_mul x332_mul_1 ( // @[Math.scala 262:24:@30183.4]
    .clock(x332_mul_1_clock),
    .io_a(x332_mul_1_io_a),
    .io_b(x332_mul_1_io_b),
    .io_flow(x332_mul_1_io_flow),
    .io_result(x332_mul_1_io_result)
  );
  x324 x333_1 ( // @[Math.scala 720:24:@30193.4]
    .io_b(x333_1_io_b),
    .io_result(x333_1_io_result)
  );
  RetimeWrapper_198 RetimeWrapper_77 ( // @[package.scala 93:22:@30202.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x314_x13 x334_sum_1 ( // @[Math.scala 150:24:@30211.4]
    .clock(x334_sum_1_clock),
    .reset(x334_sum_1_reset),
    .io_a(x334_sum_1_io_a),
    .io_b(x334_sum_1_io_b),
    .io_flow(x334_sum_1_io_flow),
    .io_result(x334_sum_1_io_result)
  );
  RetimeWrapper_286 RetimeWrapper_78 ( // @[package.scala 93:22:@30225.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_79 ( // @[package.scala 93:22:@30234.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_80 ( // @[package.scala 93:22:@30243.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_81 ( // @[package.scala 93:22:@30252.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  assign b223 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 62:18:@27791.4]
  assign b224 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 63:18:@27792.4]
  assign _T_205 = b223 & b224; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 67:30:@27794.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 67:37:@27795.4]
  assign _T_210 = io_in_x194_TID == 8'h0; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 69:76:@27800.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 69:62:@27801.4]
  assign _T_213 = io_in_x194_TDEST == 8'h0; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 69:101:@27802.4]
  assign b221_number = __io_result; // @[Math.scala 723:22:@27776.4 Math.scala 724:14:@27777.4]
  assign _T_241 = $signed(b221_number); // @[Math.scala 406:49:@27892.4]
  assign _T_243 = $signed(_T_241) & $signed(32'sh3); // @[Math.scala 406:56:@27894.4]
  assign _T_244 = $signed(_T_243); // @[Math.scala 406:56:@27895.4]
  assign x394_number = $unsigned(_T_244); // @[implicits.scala 133:21:@27896.4]
  assign _T_254 = $signed(x394_number); // @[Math.scala 406:49:@27905.4]
  assign _T_256 = $signed(_T_254) & $signed(32'sh3); // @[Math.scala 406:56:@27907.4]
  assign _T_257 = $signed(_T_256); // @[Math.scala 406:56:@27908.4]
  assign b222_number = __1_io_result; // @[Math.scala 723:22:@27788.4 Math.scala 724:14:@27789.4]
  assign _T_261 = b222_number[31]; // @[FixedPoint.scala 50:25:@27914.4]
  assign _T_265 = _T_261 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@27916.4]
  assign _T_266 = b222_number[31:16]; // @[FixedPoint.scala 18:52:@27917.4]
  assign _T_272 = _T_266 == 16'hffff; // @[Math.scala 451:55:@27919.4]
  assign _T_273 = b222_number[15:0]; // @[FixedPoint.scala 18:52:@27920.4]
  assign _T_279 = _T_273 != 16'h0; // @[Math.scala 451:110:@27922.4]
  assign _T_280 = _T_272 & _T_279; // @[Math.scala 451:94:@27923.4]
  assign _T_282 = {_T_265,_T_266}; // @[Cat.scala 30:58:@27925.4]
  assign _T_292 = $signed(b222_number); // @[Math.scala 406:49:@27933.4]
  assign _T_294 = $signed(_T_292) & $signed(32'shffff); // @[Math.scala 406:56:@27935.4]
  assign _T_295 = $signed(_T_294); // @[Math.scala 406:56:@27936.4]
  assign x398_sum_number = x398_sum_1_io_result; // @[Math.scala 154:22:@27947.4 Math.scala 155:14:@27948.4]
  assign _T_302 = x398_sum_number[31]; // @[FixedPoint.scala 50:25:@27952.4]
  assign _T_306 = _T_302 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@27954.4]
  assign _T_307 = x398_sum_number[31:8]; // @[FixedPoint.scala 18:52:@27955.4]
  assign _T_313 = _T_307 == 24'hffffff; // @[Math.scala 451:55:@27957.4]
  assign _T_314 = x398_sum_number[7:0]; // @[FixedPoint.scala 18:52:@27958.4]
  assign _T_320 = _T_314 != 8'h0; // @[Math.scala 451:110:@27960.4]
  assign _T_321 = _T_313 & _T_320; // @[Math.scala 451:94:@27961.4]
  assign _T_323 = {_T_306,_T_307}; // @[Cat.scala 30:58:@27963.4]
  assign _T_333 = $signed(x398_sum_number); // @[Math.scala 406:49:@27971.4]
  assign _T_335 = $signed(_T_333) & $signed(32'shff); // @[Math.scala 406:56:@27973.4]
  assign _T_336 = $signed(_T_335); // @[Math.scala 406:56:@27974.4]
  assign x401_sum_number = x401_sum_1_io_result; // @[Math.scala 154:22:@27985.4 Math.scala 155:14:@27986.4]
  assign _T_343 = x401_sum_number[31]; // @[FixedPoint.scala 50:25:@27990.4]
  assign _T_347 = _T_343 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@27992.4]
  assign _T_348 = x401_sum_number[31:4]; // @[FixedPoint.scala 18:52:@27993.4]
  assign _T_354 = _T_348 == 28'hfffffff; // @[Math.scala 451:55:@27995.4]
  assign _T_355 = x401_sum_number[3:0]; // @[FixedPoint.scala 18:52:@27996.4]
  assign _T_361 = _T_355 != 4'h0; // @[Math.scala 451:110:@27998.4]
  assign _T_362 = _T_354 & _T_361; // @[Math.scala 451:94:@27999.4]
  assign _T_364 = {_T_347,_T_348}; // @[Cat.scala 30:58:@28001.4]
  assign _T_374 = $signed(x401_sum_number); // @[Math.scala 406:49:@28009.4]
  assign _T_376 = $signed(_T_374) & $signed(32'shf); // @[Math.scala 406:56:@28011.4]
  assign _T_377 = $signed(_T_376); // @[Math.scala 406:56:@28012.4]
  assign x404_sum_number = x404_sum_1_io_result; // @[Math.scala 154:22:@28023.4 Math.scala 155:14:@28024.4]
  assign _T_384 = x404_sum_number[31]; // @[FixedPoint.scala 50:25:@28028.4]
  assign _T_388 = _T_384 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28030.4]
  assign _T_389 = x404_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28031.4]
  assign _T_395 = _T_389 == 30'h3fffffff; // @[Math.scala 451:55:@28033.4]
  assign _T_396 = x404_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28034.4]
  assign _T_402 = _T_396 != 2'h0; // @[Math.scala 451:110:@28036.4]
  assign _T_403 = _T_395 & _T_402; // @[Math.scala 451:94:@28037.4]
  assign _T_405 = {_T_388,_T_389}; // @[Cat.scala 30:58:@28039.4]
  assign _T_415 = $signed(x404_sum_number); // @[Math.scala 406:49:@28047.4]
  assign _T_417 = $signed(_T_415) & $signed(32'sh3); // @[Math.scala 406:56:@28049.4]
  assign _T_418 = $signed(_T_417); // @[Math.scala 406:56:@28050.4]
  assign x407_sum_number = x407_sum_1_io_result; // @[Math.scala 154:22:@28061.4 Math.scala 155:14:@28062.4]
  assign _T_425 = x407_sum_number[31]; // @[FixedPoint.scala 50:25:@28066.4]
  assign _T_429 = _T_425 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28068.4]
  assign _T_430 = x407_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28069.4]
  assign _T_436 = _T_430 == 30'h3fffffff; // @[Math.scala 451:55:@28071.4]
  assign _T_437 = x407_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28072.4]
  assign _T_443 = _T_437 != 2'h0; // @[Math.scala 451:110:@28074.4]
  assign _T_444 = _T_436 & _T_443; // @[Math.scala 451:94:@28075.4]
  assign _T_448 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@28083.4 package.scala 96:25:@28084.4]
  assign _T_458 = $signed(x407_sum_number); // @[Math.scala 406:49:@28092.4]
  assign _T_460 = $signed(_T_458) & $signed(32'sh3); // @[Math.scala 406:56:@28094.4]
  assign _T_461 = $signed(_T_460); // @[Math.scala 406:56:@28095.4]
  assign _T_465 = $signed(RetimeWrapper_2_io_out); // @[package.scala 96:25:@28103.4]
  assign x410_sum_number = x410_sum_1_io_result; // @[Math.scala 154:22:@28115.4 Math.scala 155:14:@28116.4]
  assign _T_472 = x410_sum_number[31]; // @[FixedPoint.scala 50:25:@28120.4]
  assign _T_476 = _T_472 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28122.4]
  assign _T_477 = x410_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28123.4]
  assign _T_483 = _T_477 == 30'h3fffffff; // @[Math.scala 451:55:@28125.4]
  assign _T_484 = x410_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28126.4]
  assign _T_490 = _T_484 != 2'h0; // @[Math.scala 451:110:@28128.4]
  assign _T_491 = _T_483 & _T_490; // @[Math.scala 451:94:@28129.4]
  assign _T_493 = {_T_476,_T_477}; // @[Cat.scala 30:58:@28131.4]
  assign _T_503 = $signed(x410_sum_number); // @[Math.scala 406:49:@28139.4]
  assign _T_505 = $signed(_T_503) & $signed(32'sh3); // @[Math.scala 406:56:@28141.4]
  assign _T_506 = $signed(_T_505); // @[Math.scala 406:56:@28142.4]
  assign x413_sum_number = x413_sum_1_io_result; // @[Math.scala 154:22:@28153.4 Math.scala 155:14:@28154.4]
  assign _T_516 = $signed(x413_sum_number); // @[Math.scala 476:37:@28159.4]
  assign x482_x414_D1 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@28197.4 package.scala 96:25:@28198.4]
  assign x483_x413_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@28206.4 package.scala 96:25:@28207.4]
  assign x416_sub_number = x416_sub_1_io_result; // @[Math.scala 195:22:@28179.4 Math.scala 196:14:@28180.4]
  assign _T_547 = x394_number[31]; // @[FixedPoint.scala 50:25:@28214.4]
  assign _T_551 = _T_547 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28216.4]
  assign _T_552 = x394_number[31:2]; // @[FixedPoint.scala 18:52:@28217.4]
  assign _T_558 = _T_552 == 30'h3fffffff; // @[Math.scala 451:55:@28219.4]
  assign _T_559 = x394_number[1:0]; // @[FixedPoint.scala 18:52:@28220.4]
  assign _T_565 = _T_559 != 2'h0; // @[Math.scala 451:110:@28222.4]
  assign _T_566 = _T_558 & _T_565; // @[Math.scala 451:94:@28223.4]
  assign _T_568 = {_T_551,_T_552}; // @[Cat.scala 30:58:@28225.4]
  assign x233_1_number = _T_566 ? 32'h0 : _T_568; // @[Math.scala 454:20:@28226.4]
  assign _GEN_0 = {{9'd0}, x233_1_number}; // @[Math.scala 461:32:@28231.4]
  assign _T_573 = _GEN_0 << 9; // @[Math.scala 461:32:@28231.4]
  assign _GEN_1 = {{7'd0}, x233_1_number}; // @[Math.scala 461:32:@28236.4]
  assign _T_576 = _GEN_1 << 7; // @[Math.scala 461:32:@28236.4]
  assign _T_609 = ~ io_sigsIn_break; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:101:@28325.4]
  assign _T_613 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@28333.4 package.scala 96:25:@28334.4]
  assign _T_615 = io_rr ? _T_613 : 1'h0; // @[implicits.scala 55:10:@28335.4]
  assign _T_616 = _T_609 & _T_615; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:118:@28336.4]
  assign _T_618 = _T_616 & _T_609; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:207:@28338.4]
  assign _T_619 = _T_618 & io_sigsIn_backpressure; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:226:@28339.4]
  assign x488_b223_D21 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@28313.4 package.scala 96:25:@28314.4]
  assign _T_620 = _T_619 & x488_b223_D21; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 163:252:@28340.4]
  assign x486_b224_D21 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@28295.4 package.scala 96:25:@28296.4]
  assign x490_b221_D23_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@28354.4 package.scala 96:25:@28355.4]
  assign _T_630 = $signed(x490_b221_D23_number); // @[Math.scala 476:37:@28360.4]
  assign x491_b222_D23_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@28377.4 package.scala 96:25:@28378.4]
  assign _T_645 = $signed(x491_b222_D23_number); // @[Math.scala 476:37:@28385.4]
  assign x239 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@28368.4 package.scala 96:25:@28369.4]
  assign x240 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@28393.4 package.scala 96:25:@28394.4]
  assign x241 = x239 | x240; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 182:59:@28397.4]
  assign _T_683 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@28465.4 package.scala 96:25:@28466.4]
  assign _T_685 = io_rr ? _T_683 : 1'h0; // @[implicits.scala 55:10:@28467.4]
  assign _T_686 = _T_609 & _T_685; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 201:194:@28468.4]
  assign x496_x242_D21 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@28444.4 package.scala 96:25:@28445.4]
  assign _T_687 = _T_686 & x496_x242_D21; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 201:283:@28469.4]
  assign x495_b223_D45 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@28435.4 package.scala 96:25:@28436.4]
  assign _T_688 = _T_687 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 201:291:@28470.4]
  assign x493_b224_D45 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@28417.4 package.scala 96:25:@28418.4]
  assign x245_rdcol_number = x245_rdcol_1_io_result; // @[Math.scala 195:22:@28489.4 Math.scala 196:14:@28490.4]
  assign _T_703 = $signed(x245_rdcol_number); // @[Math.scala 476:37:@28495.4]
  assign x498_x239_D1 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@28512.4 package.scala 96:25:@28513.4]
  assign x246 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@28503.4 package.scala 96:25:@28504.4]
  assign x247 = x498_x239_D1 | x246; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 211:24:@28516.4]
  assign _T_717 = x245_rdcol_number[31]; // @[FixedPoint.scala 50:25:@28523.4]
  assign _T_721 = _T_717 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@28525.4]
  assign _T_722 = x245_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@28526.4]
  assign _T_728 = _T_722 == 16'hffff; // @[Math.scala 451:55:@28528.4]
  assign _T_729 = x245_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@28529.4]
  assign _T_735 = _T_729 != 16'h0; // @[Math.scala 451:110:@28531.4]
  assign _T_736 = _T_728 & _T_735; // @[Math.scala 451:94:@28532.4]
  assign _T_738 = {_T_721,_T_722}; // @[Cat.scala 30:58:@28534.4]
  assign _T_750 = $signed(_T_703) & $signed(32'shffff); // @[Math.scala 406:56:@28544.4]
  assign _T_751 = $signed(_T_750); // @[Math.scala 406:56:@28545.4]
  assign x423_sum_number = x423_sum_1_io_result; // @[Math.scala 154:22:@28556.4 Math.scala 155:14:@28557.4]
  assign _T_758 = x423_sum_number[31]; // @[FixedPoint.scala 50:25:@28561.4]
  assign _T_762 = _T_758 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@28563.4]
  assign _T_763 = x423_sum_number[31:8]; // @[FixedPoint.scala 18:52:@28564.4]
  assign _T_769 = _T_763 == 24'hffffff; // @[Math.scala 451:55:@28566.4]
  assign _T_770 = x423_sum_number[7:0]; // @[FixedPoint.scala 18:52:@28567.4]
  assign _T_776 = _T_770 != 8'h0; // @[Math.scala 451:110:@28569.4]
  assign _T_777 = _T_769 & _T_776; // @[Math.scala 451:94:@28570.4]
  assign _T_781 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@28578.4 package.scala 96:25:@28579.4]
  assign _T_791 = $signed(x423_sum_number); // @[Math.scala 406:49:@28587.4]
  assign _T_793 = $signed(_T_791) & $signed(32'shff); // @[Math.scala 406:56:@28589.4]
  assign _T_794 = $signed(_T_793); // @[Math.scala 406:56:@28590.4]
  assign _T_798 = $signed(RetimeWrapper_27_io_out); // @[package.scala 96:25:@28598.4]
  assign x426_sum_number = x426_sum_1_io_result; // @[Math.scala 154:22:@28610.4 Math.scala 155:14:@28611.4]
  assign _T_805 = x426_sum_number[31]; // @[FixedPoint.scala 50:25:@28615.4]
  assign _T_809 = _T_805 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@28617.4]
  assign _T_810 = x426_sum_number[31:4]; // @[FixedPoint.scala 18:52:@28618.4]
  assign _T_816 = _T_810 == 28'hfffffff; // @[Math.scala 451:55:@28620.4]
  assign _T_817 = x426_sum_number[3:0]; // @[FixedPoint.scala 18:52:@28621.4]
  assign _T_823 = _T_817 != 4'h0; // @[Math.scala 451:110:@28623.4]
  assign _T_824 = _T_816 & _T_823; // @[Math.scala 451:94:@28624.4]
  assign _T_826 = {_T_809,_T_810}; // @[Cat.scala 30:58:@28626.4]
  assign _T_836 = $signed(x426_sum_number); // @[Math.scala 406:49:@28634.4]
  assign _T_838 = $signed(_T_836) & $signed(32'shf); // @[Math.scala 406:56:@28636.4]
  assign _T_839 = $signed(_T_838); // @[Math.scala 406:56:@28637.4]
  assign x429_sum_number = x429_sum_1_io_result; // @[Math.scala 154:22:@28648.4 Math.scala 155:14:@28649.4]
  assign _T_846 = x429_sum_number[31]; // @[FixedPoint.scala 50:25:@28653.4]
  assign _T_850 = _T_846 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28655.4]
  assign _T_851 = x429_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28656.4]
  assign _T_857 = _T_851 == 30'h3fffffff; // @[Math.scala 451:55:@28658.4]
  assign _T_858 = x429_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28659.4]
  assign _T_864 = _T_858 != 2'h0; // @[Math.scala 451:110:@28661.4]
  assign _T_865 = _T_857 & _T_864; // @[Math.scala 451:94:@28662.4]
  assign _T_867 = {_T_850,_T_851}; // @[Cat.scala 30:58:@28664.4]
  assign _T_877 = $signed(x429_sum_number); // @[Math.scala 406:49:@28672.4]
  assign _T_879 = $signed(_T_877) & $signed(32'sh3); // @[Math.scala 406:56:@28674.4]
  assign _T_880 = $signed(_T_879); // @[Math.scala 406:56:@28675.4]
  assign x432_sum_number = x432_sum_1_io_result; // @[Math.scala 154:22:@28686.4 Math.scala 155:14:@28687.4]
  assign _T_887 = x432_sum_number[31]; // @[FixedPoint.scala 50:25:@28691.4]
  assign _T_891 = _T_887 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28693.4]
  assign _T_892 = x432_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28694.4]
  assign _T_898 = _T_892 == 30'h3fffffff; // @[Math.scala 451:55:@28696.4]
  assign _T_899 = x432_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28697.4]
  assign _T_905 = _T_899 != 2'h0; // @[Math.scala 451:110:@28699.4]
  assign _T_906 = _T_898 & _T_905; // @[Math.scala 451:94:@28700.4]
  assign _T_908 = {_T_891,_T_892}; // @[Cat.scala 30:58:@28702.4]
  assign _T_918 = $signed(x432_sum_number); // @[Math.scala 406:49:@28710.4]
  assign _T_920 = $signed(_T_918) & $signed(32'sh3); // @[Math.scala 406:56:@28712.4]
  assign _T_921 = $signed(_T_920); // @[Math.scala 406:56:@28713.4]
  assign x435_sum_number = x435_sum_1_io_result; // @[Math.scala 154:22:@28724.4 Math.scala 155:14:@28725.4]
  assign _T_928 = x435_sum_number[31]; // @[FixedPoint.scala 50:25:@28729.4]
  assign _T_932 = _T_928 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28731.4]
  assign _T_933 = x435_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28732.4]
  assign _T_939 = _T_933 == 30'h3fffffff; // @[Math.scala 451:55:@28734.4]
  assign _T_940 = x435_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28735.4]
  assign _T_946 = _T_940 != 2'h0; // @[Math.scala 451:110:@28737.4]
  assign _T_947 = _T_939 & _T_946; // @[Math.scala 451:94:@28738.4]
  assign _T_949 = {_T_932,_T_933}; // @[Cat.scala 30:58:@28740.4]
  assign _T_959 = $signed(x435_sum_number); // @[Math.scala 406:49:@28748.4]
  assign _T_961 = $signed(_T_959) & $signed(32'sh3); // @[Math.scala 406:56:@28750.4]
  assign _T_962 = $signed(_T_961); // @[Math.scala 406:56:@28751.4]
  assign x438_sum_number = x438_sum_1_io_result; // @[Math.scala 154:22:@28762.4 Math.scala 155:14:@28763.4]
  assign _T_972 = $signed(x438_sum_number); // @[Math.scala 476:37:@28768.4]
  assign x439 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@28776.4 package.scala 96:25:@28777.4]
  assign x499_x438_sum_D1_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@28811.4 package.scala 96:25:@28812.4]
  assign x441_sub_number = x441_sub_1_io_result; // @[Math.scala 195:22:@28802.4 Math.scala 196:14:@28803.4]
  assign _T_1029 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@28875.4 package.scala 96:25:@28876.4]
  assign _T_1031 = io_rr ? _T_1029 : 1'h0; // @[implicits.scala 55:10:@28877.4]
  assign _T_1032 = _T_609 & _T_1031; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 274:194:@28878.4]
  assign x501_x248_D20 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@28854.4 package.scala 96:25:@28855.4]
  assign _T_1033 = _T_1032 & x501_x248_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 274:283:@28879.4]
  assign _T_1034 = _T_1033 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 274:291:@28880.4]
  assign x254_rdcol_number = x254_rdcol_1_io_result; // @[Math.scala 195:22:@28899.4 Math.scala 196:14:@28900.4]
  assign _T_1049 = $signed(x254_rdcol_number); // @[Math.scala 476:37:@28905.4]
  assign x255 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@28913.4 package.scala 96:25:@28914.4]
  assign x256 = x498_x239_D1 | x255; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 288:59:@28917.4]
  assign _T_1062 = x254_rdcol_number[31]; // @[FixedPoint.scala 50:25:@28926.4]
  assign _T_1066 = _T_1062 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@28928.4]
  assign _T_1067 = x254_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@28929.4]
  assign _T_1073 = _T_1067 == 16'hffff; // @[Math.scala 451:55:@28931.4]
  assign _T_1074 = x254_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@28932.4]
  assign _T_1080 = _T_1074 != 16'h0; // @[Math.scala 451:110:@28934.4]
  assign _T_1081 = _T_1073 & _T_1080; // @[Math.scala 451:94:@28935.4]
  assign _T_1083 = {_T_1066,_T_1067}; // @[Cat.scala 30:58:@28937.4]
  assign _T_1095 = $signed(_T_1049) & $signed(32'shffff); // @[Math.scala 406:56:@28947.4]
  assign _T_1096 = $signed(_T_1095); // @[Math.scala 406:56:@28948.4]
  assign x445_sum_number = x445_sum_1_io_result; // @[Math.scala 154:22:@28959.4 Math.scala 155:14:@28960.4]
  assign _T_1103 = x445_sum_number[31]; // @[FixedPoint.scala 50:25:@28964.4]
  assign _T_1107 = _T_1103 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@28966.4]
  assign _T_1108 = x445_sum_number[31:8]; // @[FixedPoint.scala 18:52:@28967.4]
  assign _T_1114 = _T_1108 == 24'hffffff; // @[Math.scala 451:55:@28969.4]
  assign _T_1115 = x445_sum_number[7:0]; // @[FixedPoint.scala 18:52:@28970.4]
  assign _T_1121 = _T_1115 != 8'h0; // @[Math.scala 451:110:@28972.4]
  assign _T_1122 = _T_1114 & _T_1121; // @[Math.scala 451:94:@28973.4]
  assign _T_1126 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@28981.4 package.scala 96:25:@28982.4]
  assign _T_1136 = $signed(x445_sum_number); // @[Math.scala 406:49:@28990.4]
  assign _T_1138 = $signed(_T_1136) & $signed(32'shff); // @[Math.scala 406:56:@28992.4]
  assign _T_1139 = $signed(_T_1138); // @[Math.scala 406:56:@28993.4]
  assign _T_1143 = $signed(RetimeWrapper_37_io_out); // @[package.scala 96:25:@29001.4]
  assign x448_sum_number = x448_sum_1_io_result; // @[Math.scala 154:22:@29013.4 Math.scala 155:14:@29014.4]
  assign _T_1150 = x448_sum_number[31]; // @[FixedPoint.scala 50:25:@29018.4]
  assign _T_1154 = _T_1150 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@29020.4]
  assign _T_1155 = x448_sum_number[31:4]; // @[FixedPoint.scala 18:52:@29021.4]
  assign _T_1161 = _T_1155 == 28'hfffffff; // @[Math.scala 451:55:@29023.4]
  assign _T_1162 = x448_sum_number[3:0]; // @[FixedPoint.scala 18:52:@29024.4]
  assign _T_1168 = _T_1162 != 4'h0; // @[Math.scala 451:110:@29026.4]
  assign _T_1169 = _T_1161 & _T_1168; // @[Math.scala 451:94:@29027.4]
  assign _T_1171 = {_T_1154,_T_1155}; // @[Cat.scala 30:58:@29029.4]
  assign _T_1181 = $signed(x448_sum_number); // @[Math.scala 406:49:@29037.4]
  assign _T_1183 = $signed(_T_1181) & $signed(32'shf); // @[Math.scala 406:56:@29039.4]
  assign _T_1184 = $signed(_T_1183); // @[Math.scala 406:56:@29040.4]
  assign x451_sum_number = x451_sum_1_io_result; // @[Math.scala 154:22:@29051.4 Math.scala 155:14:@29052.4]
  assign _T_1191 = x451_sum_number[31]; // @[FixedPoint.scala 50:25:@29056.4]
  assign _T_1195 = _T_1191 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@29058.4]
  assign _T_1196 = x451_sum_number[31:2]; // @[FixedPoint.scala 18:52:@29059.4]
  assign _T_1202 = _T_1196 == 30'h3fffffff; // @[Math.scala 451:55:@29061.4]
  assign _T_1203 = x451_sum_number[1:0]; // @[FixedPoint.scala 18:52:@29062.4]
  assign _T_1209 = _T_1203 != 2'h0; // @[Math.scala 451:110:@29064.4]
  assign _T_1210 = _T_1202 & _T_1209; // @[Math.scala 451:94:@29065.4]
  assign _T_1212 = {_T_1195,_T_1196}; // @[Cat.scala 30:58:@29067.4]
  assign _T_1222 = $signed(x451_sum_number); // @[Math.scala 406:49:@29075.4]
  assign _T_1224 = $signed(_T_1222) & $signed(32'sh3); // @[Math.scala 406:56:@29077.4]
  assign _T_1225 = $signed(_T_1224); // @[Math.scala 406:56:@29078.4]
  assign x454_sum_number = x454_sum_1_io_result; // @[Math.scala 154:22:@29089.4 Math.scala 155:14:@29090.4]
  assign _T_1232 = x454_sum_number[31]; // @[FixedPoint.scala 50:25:@29094.4]
  assign _T_1236 = _T_1232 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@29096.4]
  assign _T_1237 = x454_sum_number[31:2]; // @[FixedPoint.scala 18:52:@29097.4]
  assign _T_1243 = _T_1237 == 30'h3fffffff; // @[Math.scala 451:55:@29099.4]
  assign _T_1244 = x454_sum_number[1:0]; // @[FixedPoint.scala 18:52:@29100.4]
  assign _T_1250 = _T_1244 != 2'h0; // @[Math.scala 451:110:@29102.4]
  assign _T_1251 = _T_1243 & _T_1250; // @[Math.scala 451:94:@29103.4]
  assign _T_1253 = {_T_1236,_T_1237}; // @[Cat.scala 30:58:@29105.4]
  assign _T_1263 = $signed(x454_sum_number); // @[Math.scala 406:49:@29113.4]
  assign _T_1265 = $signed(_T_1263) & $signed(32'sh3); // @[Math.scala 406:56:@29115.4]
  assign _T_1266 = $signed(_T_1265); // @[Math.scala 406:56:@29116.4]
  assign x457_sum_number = x457_sum_1_io_result; // @[Math.scala 154:22:@29127.4 Math.scala 155:14:@29128.4]
  assign _T_1273 = x457_sum_number[31]; // @[FixedPoint.scala 50:25:@29132.4]
  assign _T_1277 = _T_1273 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@29134.4]
  assign _T_1278 = x457_sum_number[31:2]; // @[FixedPoint.scala 18:52:@29135.4]
  assign _T_1284 = _T_1278 == 30'h3fffffff; // @[Math.scala 451:55:@29137.4]
  assign _T_1285 = x457_sum_number[1:0]; // @[FixedPoint.scala 18:52:@29138.4]
  assign _T_1291 = _T_1285 != 2'h0; // @[Math.scala 451:110:@29140.4]
  assign _T_1292 = _T_1284 & _T_1291; // @[Math.scala 451:94:@29141.4]
  assign _T_1294 = {_T_1277,_T_1278}; // @[Cat.scala 30:58:@29143.4]
  assign _T_1304 = $signed(x457_sum_number); // @[Math.scala 406:49:@29151.4]
  assign _T_1306 = $signed(_T_1304) & $signed(32'sh3); // @[Math.scala 406:56:@29153.4]
  assign _T_1307 = $signed(_T_1306); // @[Math.scala 406:56:@29154.4]
  assign x460_sum_number = x460_sum_1_io_result; // @[Math.scala 154:22:@29165.4 Math.scala 155:14:@29166.4]
  assign _T_1317 = $signed(x460_sum_number); // @[Math.scala 476:37:@29171.4]
  assign x461 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@29179.4 package.scala 96:25:@29180.4]
  assign x503_x460_sum_D1_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@29214.4 package.scala 96:25:@29215.4]
  assign x463_sub_number = x463_sub_1_io_result; // @[Math.scala 195:22:@29205.4 Math.scala 196:14:@29206.4]
  assign _T_1371 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@29269.4 package.scala 96:25:@29270.4]
  assign _T_1373 = io_rr ? _T_1371 : 1'h0; // @[implicits.scala 55:10:@29271.4]
  assign _T_1374 = _T_609 & _T_1373; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 351:194:@29272.4]
  assign x504_x257_D20 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@29248.4 package.scala 96:25:@29249.4]
  assign _T_1375 = _T_1374 & x504_x257_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 351:283:@29273.4]
  assign _T_1376 = _T_1375 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 351:291:@29274.4]
  assign x263_rdrow_number = x263_rdrow_1_io_result; // @[Math.scala 195:22:@29293.4 Math.scala 196:14:@29294.4]
  assign _T_1393 = $signed(x263_rdrow_number); // @[Math.scala 406:49:@29300.4]
  assign _T_1395 = $signed(_T_1393) & $signed(32'sh3); // @[Math.scala 406:56:@29302.4]
  assign _T_1396 = $signed(_T_1395); // @[Math.scala 406:56:@29303.4]
  assign x465_number = $unsigned(_T_1396); // @[implicits.scala 133:21:@29304.4]
  assign x265 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@29318.4 package.scala 96:25:@29319.4]
  assign x506_x240_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@29327.4 package.scala 96:25:@29328.4]
  assign x266 = x265 | x506_x240_D1; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 363:24:@29331.4]
  assign _T_1422 = $signed(x465_number); // @[Math.scala 406:49:@29340.4]
  assign _T_1424 = $signed(_T_1422) & $signed(32'sh3); // @[Math.scala 406:56:@29342.4]
  assign _T_1425 = $signed(_T_1424); // @[Math.scala 406:56:@29343.4]
  assign _T_1429 = $signed(RetimeWrapper_46_io_out); // @[package.scala 96:25:@29351.4]
  assign _T_1433 = x465_number[31]; // @[FixedPoint.scala 50:25:@29358.4]
  assign _T_1437 = _T_1433 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@29360.4]
  assign _T_1438 = x465_number[31:2]; // @[FixedPoint.scala 18:52:@29361.4]
  assign _T_1444 = _T_1438 == 30'h3fffffff; // @[Math.scala 451:55:@29363.4]
  assign _T_1445 = x465_number[1:0]; // @[FixedPoint.scala 18:52:@29364.4]
  assign _T_1451 = _T_1445 != 2'h0; // @[Math.scala 451:110:@29366.4]
  assign _T_1452 = _T_1444 & _T_1451; // @[Math.scala 451:94:@29367.4]
  assign _T_1456 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@29375.4 package.scala 96:25:@29376.4]
  assign x269_1_number = _T_1452 ? 32'h0 : _T_1456; // @[Math.scala 454:20:@29377.4]
  assign _GEN_2 = {{9'd0}, x269_1_number}; // @[Math.scala 461:32:@29382.4]
  assign _T_1461 = _GEN_2 << 9; // @[Math.scala 461:32:@29382.4]
  assign _GEN_3 = {{7'd0}, x269_1_number}; // @[Math.scala 461:32:@29387.4]
  assign _T_1464 = _GEN_3 << 7; // @[Math.scala 461:32:@29387.4]
  assign _T_1497 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@29464.4 package.scala 96:25:@29465.4]
  assign _T_1499 = io_rr ? _T_1497 : 1'h0; // @[implicits.scala 55:10:@29466.4]
  assign _T_1500 = _T_609 & _T_1499; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 392:194:@29467.4]
  assign x511_x267_D20 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@29452.4 package.scala 96:25:@29453.4]
  assign _T_1501 = _T_1500 & x511_x267_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 392:283:@29468.4]
  assign _T_1502 = _T_1501 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 392:291:@29469.4]
  assign x274 = x265 | x246; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 402:59:@29480.4]
  assign _T_1531 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@29524.4 package.scala 96:25:@29525.4]
  assign _T_1533 = io_rr ? _T_1531 : 1'h0; // @[implicits.scala 55:10:@29526.4]
  assign _T_1534 = _T_609 & _T_1533; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 417:194:@29527.4]
  assign x513_x275_D20 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@29512.4 package.scala 96:25:@29513.4]
  assign _T_1535 = _T_1534 & x513_x275_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 417:283:@29528.4]
  assign _T_1536 = _T_1535 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 417:291:@29529.4]
  assign x279 = x265 | x255; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 421:59:@29540.4]
  assign _T_1560 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@29573.4 package.scala 96:25:@29574.4]
  assign _T_1562 = io_rr ? _T_1560 : 1'h0; // @[implicits.scala 55:10:@29575.4]
  assign _T_1563 = _T_609 & _T_1562; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 432:194:@29576.4]
  assign x514_x280_D20 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@29561.4 package.scala 96:25:@29562.4]
  assign _T_1564 = _T_1563 & x514_x280_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 432:283:@29577.4]
  assign _T_1565 = _T_1564 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 432:291:@29578.4]
  assign x284_rdrow_number = x284_rdrow_1_io_result; // @[Math.scala 195:22:@29597.4 Math.scala 196:14:@29598.4]
  assign _T_1582 = $signed(x284_rdrow_number); // @[Math.scala 406:49:@29604.4]
  assign _T_1584 = $signed(_T_1582) & $signed(32'sh3); // @[Math.scala 406:56:@29606.4]
  assign _T_1585 = $signed(_T_1584); // @[Math.scala 406:56:@29607.4]
  assign x470_number = $unsigned(_T_1585); // @[implicits.scala 133:21:@29608.4]
  assign x286 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@29622.4 package.scala 96:25:@29623.4]
  assign x287 = x286 | x506_x240_D1; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 442:24:@29626.4]
  assign _T_1608 = $signed(x470_number); // @[Math.scala 406:49:@29635.4]
  assign _T_1610 = $signed(_T_1608) & $signed(32'sh3); // @[Math.scala 406:56:@29637.4]
  assign _T_1611 = $signed(_T_1610); // @[Math.scala 406:56:@29638.4]
  assign _T_1615 = $signed(RetimeWrapper_60_io_out); // @[package.scala 96:25:@29646.4]
  assign _T_1619 = x470_number[31]; // @[FixedPoint.scala 50:25:@29653.4]
  assign _T_1623 = _T_1619 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@29655.4]
  assign _T_1624 = x470_number[31:2]; // @[FixedPoint.scala 18:52:@29656.4]
  assign _T_1630 = _T_1624 == 30'h3fffffff; // @[Math.scala 451:55:@29658.4]
  assign _T_1631 = x470_number[1:0]; // @[FixedPoint.scala 18:52:@29659.4]
  assign _T_1637 = _T_1631 != 2'h0; // @[Math.scala 451:110:@29661.4]
  assign _T_1638 = _T_1630 & _T_1637; // @[Math.scala 451:94:@29662.4]
  assign _T_1642 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@29670.4 package.scala 96:25:@29671.4]
  assign x290_1_number = _T_1638 ? 32'h0 : _T_1642; // @[Math.scala 454:20:@29672.4]
  assign _GEN_4 = {{9'd0}, x290_1_number}; // @[Math.scala 461:32:@29677.4]
  assign _T_1647 = _GEN_4 << 9; // @[Math.scala 461:32:@29677.4]
  assign _GEN_5 = {{7'd0}, x290_1_number}; // @[Math.scala 461:32:@29682.4]
  assign _T_1650 = _GEN_5 << 7; // @[Math.scala 461:32:@29682.4]
  assign _T_1680 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@29750.4 package.scala 96:25:@29751.4]
  assign _T_1682 = io_rr ? _T_1680 : 1'h0; // @[implicits.scala 55:10:@29752.4]
  assign _T_1683 = _T_609 & _T_1682; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 469:194:@29753.4]
  assign x516_x288_D20 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@29720.4 package.scala 96:25:@29721.4]
  assign _T_1684 = _T_1683 & x516_x288_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 469:283:@29754.4]
  assign _T_1685 = _T_1684 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 469:291:@29755.4]
  assign x295 = x286 | x246; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 473:24:@29766.4]
  assign _T_1712 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@29808.4 package.scala 96:25:@29809.4]
  assign _T_1714 = io_rr ? _T_1712 : 1'h0; // @[implicits.scala 55:10:@29810.4]
  assign _T_1715 = _T_609 & _T_1714; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 486:194:@29811.4]
  assign x520_x296_D20 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@29796.4 package.scala 96:25:@29797.4]
  assign _T_1716 = _T_1715 & x520_x296_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 486:283:@29812.4]
  assign _T_1717 = _T_1716 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 486:291:@29813.4]
  assign x300 = x286 | x255; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 490:24:@29824.4]
  assign _T_1741 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@29857.4 package.scala 96:25:@29858.4]
  assign _T_1743 = io_rr ? _T_1741 : 1'h0; // @[implicits.scala 55:10:@29859.4]
  assign _T_1744 = _T_609 & _T_1743; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 501:194:@29860.4]
  assign x521_x301_D20 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@29845.4 package.scala 96:25:@29846.4]
  assign _T_1745 = _T_1744 & x521_x301_D20; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 501:283:@29861.4]
  assign _T_1746 = _T_1745 & x495_b223_D45; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 501:291:@29862.4]
  assign x325_sub_number = x325_sub_1_io_result; // @[Math.scala 195:22:@30117.4 Math.scala 196:14:@30118.4]
  assign x327_sub_number = x327_sub_1_io_result; // @[Math.scala 195:22:@30139.4 Math.scala 196:14:@30140.4]
  assign x326 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@30129.4 package.scala 96:25:@30130.4]
  assign x328 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@30151.4 package.scala 96:25:@30152.4]
  assign x329 = x326 | x328; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 565:24:@30155.4]
  assign x524_x325_sub_D1_number = RetimeWrapper_76_io_out; // @[package.scala 96:25:@30163.4 package.scala 96:25:@30164.4]
  assign _T_1928 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@30257.4 package.scala 96:25:@30258.4]
  assign _T_1930 = io_rr ? _T_1928 : 1'h0; // @[implicits.scala 55:10:@30259.4]
  assign x526_b223_D75 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@30239.4 package.scala 96:25:@30240.4]
  assign _T_1931 = _T_1930 & x526_b223_D75; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 589:117:@30260.4]
  assign x527_b224_D75 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@30248.4 package.scala 96:25:@30249.4]
  assign _T_1932 = _T_1931 & x527_b224_D75; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 589:123:@30261.4]
  assign x236_sum_number = x236_sum_1_io_result; // @[Math.scala 154:22:@28277.4 Math.scala 155:14:@28278.4]
  assign x485_x417_D13_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@28286.4 package.scala 96:25:@28287.4]
  assign x489_x395_D21_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@28322.4 package.scala 96:25:@28323.4]
  assign x492_x417_D37_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@28408.4 package.scala 96:25:@28409.4]
  assign x494_x236_sum_D24_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@28426.4 package.scala 96:25:@28427.4]
  assign x497_x395_D45_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@28453.4 package.scala 96:25:@28454.4]
  assign x251_sum_number = x251_sum_1_io_result; // @[Math.scala 154:22:@28845.4 Math.scala 155:14:@28846.4]
  assign x502_x442_D13_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@28863.4 package.scala 96:25:@28864.4]
  assign x260_sum_number = x260_sum_1_io_result; // @[Math.scala 154:22:@29239.4 Math.scala 155:14:@29240.4]
  assign x505_x464_D13_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@29257.4 package.scala 96:25:@29258.4]
  assign x509_x466_D20_number = RetimeWrapper_50_io_out; // @[package.scala 96:25:@29434.4 package.scala 96:25:@29435.4]
  assign x510_x271_sum_D1_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@29443.4 package.scala 96:25:@29444.4]
  assign x276_sum_number = x276_sum_1_io_result; // @[Math.scala 154:22:@29503.4 Math.scala 155:14:@29504.4]
  assign x281_sum_number = x281_sum_1_io_result; // @[Math.scala 154:22:@29552.4 Math.scala 155:14:@29553.4]
  assign x517_x292_sum_D1_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@29729.4 package.scala 96:25:@29730.4]
  assign x518_x471_D20_number = RetimeWrapper_65_io_out; // @[package.scala 96:25:@29738.4 package.scala 96:25:@29739.4]
  assign x297_sum_number = x297_sum_1_io_result; // @[Math.scala 154:22:@29787.4 Math.scala 155:14:@29788.4]
  assign x302_sum_number = x302_sum_1_io_result; // @[Math.scala 154:22:@29836.4 Math.scala 155:14:@29837.4]
  assign io_in_x194_TREADY = _T_211 & _T_213; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 67:22:@27796.4 sm_x339_inr_Foreach_SAMPLER_BOX.scala 69:22:@27804.4]
  assign io_in_x195_TVALID = _T_1932 & io_sigsIn_backpressure; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 589:22:@30263.4]
  assign io_in_x195_TDATA = {{224'd0}, RetimeWrapper_78_io_out}; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 590:24:@30264.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@27774.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@27786.4]
  assign RetimeWrapper_clock = clock; // @[:@27807.4]
  assign RetimeWrapper_reset = reset; // @[:@27808.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27810.4]
  assign RetimeWrapper_io_in = io_in_x194_TDATA[31:0]; // @[package.scala 94:16:@27809.4]
  assign x227_lb_0_clock = clock; // @[:@27817.4]
  assign x227_lb_0_reset = reset; // @[:@27818.4]
  assign x227_lb_0_io_rPort_8_banks_1 = x502_x442_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@29532.4]
  assign x227_lb_0_io_rPort_8_banks_0 = x509_x466_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29531.4]
  assign x227_lb_0_io_rPort_8_ofs_0 = x276_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29533.4]
  assign x227_lb_0_io_rPort_8_en_0 = _T_1536 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@29535.4]
  assign x227_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29534.4]
  assign x227_lb_0_io_rPort_7_banks_1 = x492_x417_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@29472.4]
  assign x227_lb_0_io_rPort_7_banks_0 = x509_x466_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29471.4]
  assign x227_lb_0_io_rPort_7_ofs_0 = x510_x271_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@29473.4]
  assign x227_lb_0_io_rPort_7_en_0 = _T_1502 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@29475.4]
  assign x227_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29474.4]
  assign x227_lb_0_io_rPort_6_banks_1 = x505_x464_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@29581.4]
  assign x227_lb_0_io_rPort_6_banks_0 = x509_x466_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29580.4]
  assign x227_lb_0_io_rPort_6_ofs_0 = x281_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29582.4]
  assign x227_lb_0_io_rPort_6_en_0 = _T_1565 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@29584.4]
  assign x227_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29583.4]
  assign x227_lb_0_io_rPort_5_banks_1 = x505_x464_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@29865.4]
  assign x227_lb_0_io_rPort_5_banks_0 = x518_x471_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29864.4]
  assign x227_lb_0_io_rPort_5_ofs_0 = x302_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29866.4]
  assign x227_lb_0_io_rPort_5_en_0 = _T_1746 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@29868.4]
  assign x227_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29867.4]
  assign x227_lb_0_io_rPort_4_banks_1 = x502_x442_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@29816.4]
  assign x227_lb_0_io_rPort_4_banks_0 = x518_x471_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29815.4]
  assign x227_lb_0_io_rPort_4_ofs_0 = x297_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29817.4]
  assign x227_lb_0_io_rPort_4_en_0 = _T_1717 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@29819.4]
  assign x227_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29818.4]
  assign x227_lb_0_io_rPort_3_banks_1 = x502_x442_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@28883.4]
  assign x227_lb_0_io_rPort_3_banks_0 = x497_x395_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@28882.4]
  assign x227_lb_0_io_rPort_3_ofs_0 = x251_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28884.4]
  assign x227_lb_0_io_rPort_3_en_0 = _T_1034 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@28886.4]
  assign x227_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28885.4]
  assign x227_lb_0_io_rPort_2_banks_1 = x492_x417_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@28473.4]
  assign x227_lb_0_io_rPort_2_banks_0 = x497_x395_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@28472.4]
  assign x227_lb_0_io_rPort_2_ofs_0 = x494_x236_sum_D24_number[9:0]; // @[MemInterfaceType.scala 107:54:@28474.4]
  assign x227_lb_0_io_rPort_2_en_0 = _T_688 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@28476.4]
  assign x227_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28475.4]
  assign x227_lb_0_io_rPort_1_banks_1 = x492_x417_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@29758.4]
  assign x227_lb_0_io_rPort_1_banks_0 = x518_x471_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29757.4]
  assign x227_lb_0_io_rPort_1_ofs_0 = x517_x292_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@29759.4]
  assign x227_lb_0_io_rPort_1_en_0 = _T_1685 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@29761.4]
  assign x227_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29760.4]
  assign x227_lb_0_io_rPort_0_banks_1 = x505_x464_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@29277.4]
  assign x227_lb_0_io_rPort_0_banks_0 = x497_x395_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@29276.4]
  assign x227_lb_0_io_rPort_0_ofs_0 = x260_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29278.4]
  assign x227_lb_0_io_rPort_0_en_0 = _T_1376 & x493_b224_D45; // @[MemInterfaceType.scala 110:79:@29280.4]
  assign x227_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29279.4]
  assign x227_lb_0_io_wPort_0_banks_1 = x485_x417_D13_number[1:0]; // @[MemInterfaceType.scala 88:58:@28343.4]
  assign x227_lb_0_io_wPort_0_banks_0 = x489_x395_D21_number[2:0]; // @[MemInterfaceType.scala 88:58:@28342.4]
  assign x227_lb_0_io_wPort_0_ofs_0 = x236_sum_number[9:0]; // @[MemInterfaceType.scala 89:54:@28344.4]
  assign x227_lb_0_io_wPort_0_data_0 = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 90:56:@28345.4]
  assign x227_lb_0_io_wPort_0_en_0 = _T_620 & x486_b224_D21; // @[MemInterfaceType.scala 93:57:@28347.4]
  assign x398_sum_1_clock = clock; // @[:@27942.4]
  assign x398_sum_1_reset = reset; // @[:@27943.4]
  assign x398_sum_1_io_a = _T_280 ? 32'h0 : _T_282; // @[Math.scala 151:17:@27944.4]
  assign x398_sum_1_io_b = $unsigned(_T_295); // @[Math.scala 152:17:@27945.4]
  assign x398_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@27946.4]
  assign x401_sum_1_clock = clock; // @[:@27980.4]
  assign x401_sum_1_reset = reset; // @[:@27981.4]
  assign x401_sum_1_io_a = _T_321 ? 32'h0 : _T_323; // @[Math.scala 151:17:@27982.4]
  assign x401_sum_1_io_b = $unsigned(_T_336); // @[Math.scala 152:17:@27983.4]
  assign x401_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@27984.4]
  assign x404_sum_1_clock = clock; // @[:@28018.4]
  assign x404_sum_1_reset = reset; // @[:@28019.4]
  assign x404_sum_1_io_a = _T_362 ? 32'h0 : _T_364; // @[Math.scala 151:17:@28020.4]
  assign x404_sum_1_io_b = $unsigned(_T_377); // @[Math.scala 152:17:@28021.4]
  assign x404_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28022.4]
  assign x407_sum_1_clock = clock; // @[:@28056.4]
  assign x407_sum_1_reset = reset; // @[:@28057.4]
  assign x407_sum_1_io_a = _T_403 ? 32'h0 : _T_405; // @[Math.scala 151:17:@28058.4]
  assign x407_sum_1_io_b = $unsigned(_T_418); // @[Math.scala 152:17:@28059.4]
  assign x407_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28060.4]
  assign RetimeWrapper_1_clock = clock; // @[:@28079.4]
  assign RetimeWrapper_1_reset = reset; // @[:@28080.4]
  assign RetimeWrapper_1_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28082.4]
  assign RetimeWrapper_1_io_in = {_T_429,_T_430}; // @[package.scala 94:16:@28081.4]
  assign RetimeWrapper_2_clock = clock; // @[:@28097.4]
  assign RetimeWrapper_2_reset = reset; // @[:@28098.4]
  assign RetimeWrapper_2_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28101.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_461); // @[package.scala 94:16:@28100.4]
  assign x410_sum_1_clock = clock; // @[:@28110.4]
  assign x410_sum_1_reset = reset; // @[:@28111.4]
  assign x410_sum_1_io_a = _T_444 ? 32'h0 : _T_448; // @[Math.scala 151:17:@28112.4]
  assign x410_sum_1_io_b = $unsigned(_T_465); // @[Math.scala 152:17:@28113.4]
  assign x410_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28114.4]
  assign x413_sum_1_clock = clock; // @[:@28148.4]
  assign x413_sum_1_reset = reset; // @[:@28149.4]
  assign x413_sum_1_io_a = _T_491 ? 32'h0 : _T_493; // @[Math.scala 151:17:@28150.4]
  assign x413_sum_1_io_b = $unsigned(_T_506); // @[Math.scala 152:17:@28151.4]
  assign x413_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28152.4]
  assign x416_sub_1_clock = clock; // @[:@28174.4]
  assign x416_sub_1_reset = reset; // @[:@28175.4]
  assign x416_sub_1_io_a = x413_sum_1_io_result; // @[Math.scala 192:17:@28176.4]
  assign x416_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@28177.4]
  assign x416_sub_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@28178.4]
  assign RetimeWrapper_3_clock = clock; // @[:@28184.4]
  assign RetimeWrapper_3_reset = reset; // @[:@28185.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28187.4]
  assign RetimeWrapper_3_io_in = $signed(_T_516) < $signed(32'sh6); // @[package.scala 94:16:@28186.4]
  assign RetimeWrapper_4_clock = clock; // @[:@28193.4]
  assign RetimeWrapper_4_reset = reset; // @[:@28194.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28196.4]
  assign RetimeWrapper_4_io_in = $signed(_T_516) < $signed(32'sh3); // @[package.scala 94:16:@28195.4]
  assign RetimeWrapper_5_clock = clock; // @[:@28202.4]
  assign RetimeWrapper_5_reset = reset; // @[:@28203.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28205.4]
  assign RetimeWrapper_5_io_in = x413_sum_1_io_result; // @[package.scala 94:16:@28204.4]
  assign x420_sum_1_clock = clock; // @[:@28241.4]
  assign x420_sum_1_reset = reset; // @[:@28242.4]
  assign x420_sum_1_io_a = _T_573[31:0]; // @[Math.scala 151:17:@28243.4]
  assign x420_sum_1_io_b = _T_576[31:0]; // @[Math.scala 152:17:@28244.4]
  assign x420_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28245.4]
  assign x235_div_1_clock = clock; // @[:@28253.4]
  assign x235_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@28255.4]
  assign x235_div_1_io_flow = io_in_x195_TREADY; // @[Math.scala 330:20:@28257.4]
  assign RetimeWrapper_6_clock = clock; // @[:@28263.4]
  assign RetimeWrapper_6_reset = reset; // @[:@28264.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28266.4]
  assign RetimeWrapper_6_io_in = x420_sum_1_io_result; // @[package.scala 94:16:@28265.4]
  assign x236_sum_1_clock = clock; // @[:@28272.4]
  assign x236_sum_1_reset = reset; // @[:@28273.4]
  assign x236_sum_1_io_a = RetimeWrapper_6_io_out; // @[Math.scala 151:17:@28274.4]
  assign x236_sum_1_io_b = x235_div_1_io_result; // @[Math.scala 152:17:@28275.4]
  assign x236_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28276.4]
  assign RetimeWrapper_7_clock = clock; // @[:@28282.4]
  assign RetimeWrapper_7_reset = reset; // @[:@28283.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28285.4]
  assign RetimeWrapper_7_io_in = x482_x414_D1 ? x483_x413_sum_D1_number : x416_sub_number; // @[package.scala 94:16:@28284.4]
  assign RetimeWrapper_8_clock = clock; // @[:@28291.4]
  assign RetimeWrapper_8_reset = reset; // @[:@28292.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28294.4]
  assign RetimeWrapper_8_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@28293.4]
  assign RetimeWrapper_9_clock = clock; // @[:@28300.4]
  assign RetimeWrapper_9_reset = reset; // @[:@28301.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28303.4]
  assign RetimeWrapper_9_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@28302.4]
  assign RetimeWrapper_10_clock = clock; // @[:@28309.4]
  assign RetimeWrapper_10_reset = reset; // @[:@28310.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28312.4]
  assign RetimeWrapper_10_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@28311.4]
  assign RetimeWrapper_11_clock = clock; // @[:@28318.4]
  assign RetimeWrapper_11_reset = reset; // @[:@28319.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28321.4]
  assign RetimeWrapper_11_io_in = $unsigned(_T_257); // @[package.scala 94:16:@28320.4]
  assign RetimeWrapper_12_clock = clock; // @[:@28329.4]
  assign RetimeWrapper_12_reset = reset; // @[:@28330.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28332.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28331.4]
  assign RetimeWrapper_13_clock = clock; // @[:@28350.4]
  assign RetimeWrapper_13_reset = reset; // @[:@28351.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28353.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@28352.4]
  assign RetimeWrapper_14_clock = clock; // @[:@28364.4]
  assign RetimeWrapper_14_reset = reset; // @[:@28365.4]
  assign RetimeWrapper_14_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28367.4]
  assign RetimeWrapper_14_io_in = $signed(_T_630) < $signed(32'sh0); // @[package.scala 94:16:@28366.4]
  assign RetimeWrapper_15_clock = clock; // @[:@28373.4]
  assign RetimeWrapper_15_reset = reset; // @[:@28374.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28376.4]
  assign RetimeWrapper_15_io_in = __1_io_result; // @[package.scala 94:16:@28375.4]
  assign RetimeWrapper_16_clock = clock; // @[:@28389.4]
  assign RetimeWrapper_16_reset = reset; // @[:@28390.4]
  assign RetimeWrapper_16_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28392.4]
  assign RetimeWrapper_16_io_in = $signed(_T_645) < $signed(32'sh0); // @[package.scala 94:16:@28391.4]
  assign RetimeWrapper_17_clock = clock; // @[:@28404.4]
  assign RetimeWrapper_17_reset = reset; // @[:@28405.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28407.4]
  assign RetimeWrapper_17_io_in = x482_x414_D1 ? x483_x413_sum_D1_number : x416_sub_number; // @[package.scala 94:16:@28406.4]
  assign RetimeWrapper_18_clock = clock; // @[:@28413.4]
  assign RetimeWrapper_18_reset = reset; // @[:@28414.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28416.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@28415.4]
  assign RetimeWrapper_19_clock = clock; // @[:@28422.4]
  assign RetimeWrapper_19_reset = reset; // @[:@28423.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28425.4]
  assign RetimeWrapper_19_io_in = x236_sum_1_io_result; // @[package.scala 94:16:@28424.4]
  assign RetimeWrapper_20_clock = clock; // @[:@28431.4]
  assign RetimeWrapper_20_reset = reset; // @[:@28432.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28434.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@28433.4]
  assign RetimeWrapper_21_clock = clock; // @[:@28440.4]
  assign RetimeWrapper_21_reset = reset; // @[:@28441.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28443.4]
  assign RetimeWrapper_21_io_in = ~ x241; // @[package.scala 94:16:@28442.4]
  assign RetimeWrapper_22_clock = clock; // @[:@28449.4]
  assign RetimeWrapper_22_reset = reset; // @[:@28450.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28452.4]
  assign RetimeWrapper_22_io_in = $unsigned(_T_257); // @[package.scala 94:16:@28451.4]
  assign RetimeWrapper_23_clock = clock; // @[:@28461.4]
  assign RetimeWrapper_23_reset = reset; // @[:@28462.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28464.4]
  assign RetimeWrapper_23_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28463.4]
  assign x245_rdcol_1_clock = clock; // @[:@28484.4]
  assign x245_rdcol_1_reset = reset; // @[:@28485.4]
  assign x245_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@28486.4]
  assign x245_rdcol_1_io_b = 32'h1; // @[Math.scala 193:17:@28487.4]
  assign x245_rdcol_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@28488.4]
  assign RetimeWrapper_24_clock = clock; // @[:@28499.4]
  assign RetimeWrapper_24_reset = reset; // @[:@28500.4]
  assign RetimeWrapper_24_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28502.4]
  assign RetimeWrapper_24_io_in = $signed(_T_703) < $signed(32'sh0); // @[package.scala 94:16:@28501.4]
  assign RetimeWrapper_25_clock = clock; // @[:@28508.4]
  assign RetimeWrapper_25_reset = reset; // @[:@28509.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28511.4]
  assign RetimeWrapper_25_io_in = RetimeWrapper_14_io_out; // @[package.scala 94:16:@28510.4]
  assign x423_sum_1_clock = clock; // @[:@28551.4]
  assign x423_sum_1_reset = reset; // @[:@28552.4]
  assign x423_sum_1_io_a = _T_736 ? 32'h0 : _T_738; // @[Math.scala 151:17:@28553.4]
  assign x423_sum_1_io_b = $unsigned(_T_751); // @[Math.scala 152:17:@28554.4]
  assign x423_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28555.4]
  assign RetimeWrapper_26_clock = clock; // @[:@28574.4]
  assign RetimeWrapper_26_reset = reset; // @[:@28575.4]
  assign RetimeWrapper_26_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28577.4]
  assign RetimeWrapper_26_io_in = {_T_762,_T_763}; // @[package.scala 94:16:@28576.4]
  assign RetimeWrapper_27_clock = clock; // @[:@28592.4]
  assign RetimeWrapper_27_reset = reset; // @[:@28593.4]
  assign RetimeWrapper_27_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28596.4]
  assign RetimeWrapper_27_io_in = $unsigned(_T_794); // @[package.scala 94:16:@28595.4]
  assign x426_sum_1_clock = clock; // @[:@28605.4]
  assign x426_sum_1_reset = reset; // @[:@28606.4]
  assign x426_sum_1_io_a = _T_777 ? 32'h0 : _T_781; // @[Math.scala 151:17:@28607.4]
  assign x426_sum_1_io_b = $unsigned(_T_798); // @[Math.scala 152:17:@28608.4]
  assign x426_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28609.4]
  assign x429_sum_1_clock = clock; // @[:@28643.4]
  assign x429_sum_1_reset = reset; // @[:@28644.4]
  assign x429_sum_1_io_a = _T_824 ? 32'h0 : _T_826; // @[Math.scala 151:17:@28645.4]
  assign x429_sum_1_io_b = $unsigned(_T_839); // @[Math.scala 152:17:@28646.4]
  assign x429_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28647.4]
  assign x432_sum_1_clock = clock; // @[:@28681.4]
  assign x432_sum_1_reset = reset; // @[:@28682.4]
  assign x432_sum_1_io_a = _T_865 ? 32'h0 : _T_867; // @[Math.scala 151:17:@28683.4]
  assign x432_sum_1_io_b = $unsigned(_T_880); // @[Math.scala 152:17:@28684.4]
  assign x432_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28685.4]
  assign x435_sum_1_clock = clock; // @[:@28719.4]
  assign x435_sum_1_reset = reset; // @[:@28720.4]
  assign x435_sum_1_io_a = _T_906 ? 32'h0 : _T_908; // @[Math.scala 151:17:@28721.4]
  assign x435_sum_1_io_b = $unsigned(_T_921); // @[Math.scala 152:17:@28722.4]
  assign x435_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28723.4]
  assign x438_sum_1_clock = clock; // @[:@28757.4]
  assign x438_sum_1_reset = reset; // @[:@28758.4]
  assign x438_sum_1_io_a = _T_947 ? 32'h0 : _T_949; // @[Math.scala 151:17:@28759.4]
  assign x438_sum_1_io_b = $unsigned(_T_962); // @[Math.scala 152:17:@28760.4]
  assign x438_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28761.4]
  assign RetimeWrapper_28_clock = clock; // @[:@28772.4]
  assign RetimeWrapper_28_reset = reset; // @[:@28773.4]
  assign RetimeWrapper_28_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28775.4]
  assign RetimeWrapper_28_io_in = $signed(_T_972) < $signed(32'sh3); // @[package.scala 94:16:@28774.4]
  assign RetimeWrapper_29_clock = clock; // @[:@28786.4]
  assign RetimeWrapper_29_reset = reset; // @[:@28787.4]
  assign RetimeWrapper_29_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28789.4]
  assign RetimeWrapper_29_io_in = $signed(_T_972) < $signed(32'sh6); // @[package.scala 94:16:@28788.4]
  assign x441_sub_1_clock = clock; // @[:@28797.4]
  assign x441_sub_1_reset = reset; // @[:@28798.4]
  assign x441_sub_1_io_a = x438_sum_1_io_result; // @[Math.scala 192:17:@28799.4]
  assign x441_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@28800.4]
  assign x441_sub_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@28801.4]
  assign RetimeWrapper_30_clock = clock; // @[:@28807.4]
  assign RetimeWrapper_30_reset = reset; // @[:@28808.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28810.4]
  assign RetimeWrapper_30_io_in = x438_sum_1_io_result; // @[package.scala 94:16:@28809.4]
  assign x250_div_1_clock = clock; // @[:@28821.4]
  assign x250_div_1_io_a = x245_rdcol_1_io_result; // @[Math.scala 328:17:@28823.4]
  assign x250_div_1_io_flow = io_in_x195_TREADY; // @[Math.scala 330:20:@28825.4]
  assign RetimeWrapper_31_clock = clock; // @[:@28831.4]
  assign RetimeWrapper_31_reset = reset; // @[:@28832.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28834.4]
  assign RetimeWrapper_31_io_in = x420_sum_1_io_result; // @[package.scala 94:16:@28833.4]
  assign x251_sum_1_clock = clock; // @[:@28840.4]
  assign x251_sum_1_reset = reset; // @[:@28841.4]
  assign x251_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@28842.4]
  assign x251_sum_1_io_b = x250_div_1_io_result; // @[Math.scala 152:17:@28843.4]
  assign x251_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28844.4]
  assign RetimeWrapper_32_clock = clock; // @[:@28850.4]
  assign RetimeWrapper_32_reset = reset; // @[:@28851.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28853.4]
  assign RetimeWrapper_32_io_in = ~ x247; // @[package.scala 94:16:@28852.4]
  assign RetimeWrapper_33_clock = clock; // @[:@28859.4]
  assign RetimeWrapper_33_reset = reset; // @[:@28860.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28862.4]
  assign RetimeWrapper_33_io_in = x439 ? x499_x438_sum_D1_number : x441_sub_number; // @[package.scala 94:16:@28861.4]
  assign RetimeWrapper_34_clock = clock; // @[:@28871.4]
  assign RetimeWrapper_34_reset = reset; // @[:@28872.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28874.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28873.4]
  assign x254_rdcol_1_clock = clock; // @[:@28894.4]
  assign x254_rdcol_1_reset = reset; // @[:@28895.4]
  assign x254_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@28896.4]
  assign x254_rdcol_1_io_b = 32'h2; // @[Math.scala 193:17:@28897.4]
  assign x254_rdcol_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@28898.4]
  assign RetimeWrapper_35_clock = clock; // @[:@28909.4]
  assign RetimeWrapper_35_reset = reset; // @[:@28910.4]
  assign RetimeWrapper_35_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28912.4]
  assign RetimeWrapper_35_io_in = $signed(_T_1049) < $signed(32'sh0); // @[package.scala 94:16:@28911.4]
  assign x445_sum_1_clock = clock; // @[:@28954.4]
  assign x445_sum_1_reset = reset; // @[:@28955.4]
  assign x445_sum_1_io_a = _T_1081 ? 32'h0 : _T_1083; // @[Math.scala 151:17:@28956.4]
  assign x445_sum_1_io_b = $unsigned(_T_1096); // @[Math.scala 152:17:@28957.4]
  assign x445_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@28958.4]
  assign RetimeWrapper_36_clock = clock; // @[:@28977.4]
  assign RetimeWrapper_36_reset = reset; // @[:@28978.4]
  assign RetimeWrapper_36_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28980.4]
  assign RetimeWrapper_36_io_in = {_T_1107,_T_1108}; // @[package.scala 94:16:@28979.4]
  assign RetimeWrapper_37_clock = clock; // @[:@28995.4]
  assign RetimeWrapper_37_reset = reset; // @[:@28996.4]
  assign RetimeWrapper_37_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@28999.4]
  assign RetimeWrapper_37_io_in = $unsigned(_T_1139); // @[package.scala 94:16:@28998.4]
  assign x448_sum_1_clock = clock; // @[:@29008.4]
  assign x448_sum_1_reset = reset; // @[:@29009.4]
  assign x448_sum_1_io_a = _T_1122 ? 32'h0 : _T_1126; // @[Math.scala 151:17:@29010.4]
  assign x448_sum_1_io_b = $unsigned(_T_1143); // @[Math.scala 152:17:@29011.4]
  assign x448_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29012.4]
  assign x451_sum_1_clock = clock; // @[:@29046.4]
  assign x451_sum_1_reset = reset; // @[:@29047.4]
  assign x451_sum_1_io_a = _T_1169 ? 32'h0 : _T_1171; // @[Math.scala 151:17:@29048.4]
  assign x451_sum_1_io_b = $unsigned(_T_1184); // @[Math.scala 152:17:@29049.4]
  assign x451_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29050.4]
  assign x454_sum_1_clock = clock; // @[:@29084.4]
  assign x454_sum_1_reset = reset; // @[:@29085.4]
  assign x454_sum_1_io_a = _T_1210 ? 32'h0 : _T_1212; // @[Math.scala 151:17:@29086.4]
  assign x454_sum_1_io_b = $unsigned(_T_1225); // @[Math.scala 152:17:@29087.4]
  assign x454_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29088.4]
  assign x457_sum_1_clock = clock; // @[:@29122.4]
  assign x457_sum_1_reset = reset; // @[:@29123.4]
  assign x457_sum_1_io_a = _T_1251 ? 32'h0 : _T_1253; // @[Math.scala 151:17:@29124.4]
  assign x457_sum_1_io_b = $unsigned(_T_1266); // @[Math.scala 152:17:@29125.4]
  assign x457_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29126.4]
  assign x460_sum_1_clock = clock; // @[:@29160.4]
  assign x460_sum_1_reset = reset; // @[:@29161.4]
  assign x460_sum_1_io_a = _T_1292 ? 32'h0 : _T_1294; // @[Math.scala 151:17:@29162.4]
  assign x460_sum_1_io_b = $unsigned(_T_1307); // @[Math.scala 152:17:@29163.4]
  assign x460_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29164.4]
  assign RetimeWrapper_38_clock = clock; // @[:@29175.4]
  assign RetimeWrapper_38_reset = reset; // @[:@29176.4]
  assign RetimeWrapper_38_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29178.4]
  assign RetimeWrapper_38_io_in = $signed(_T_1317) < $signed(32'sh3); // @[package.scala 94:16:@29177.4]
  assign RetimeWrapper_39_clock = clock; // @[:@29189.4]
  assign RetimeWrapper_39_reset = reset; // @[:@29190.4]
  assign RetimeWrapper_39_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29192.4]
  assign RetimeWrapper_39_io_in = $signed(_T_1317) < $signed(32'sh6); // @[package.scala 94:16:@29191.4]
  assign x463_sub_1_clock = clock; // @[:@29200.4]
  assign x463_sub_1_reset = reset; // @[:@29201.4]
  assign x463_sub_1_io_a = x460_sum_1_io_result; // @[Math.scala 192:17:@29202.4]
  assign x463_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@29203.4]
  assign x463_sub_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@29204.4]
  assign RetimeWrapper_40_clock = clock; // @[:@29210.4]
  assign RetimeWrapper_40_reset = reset; // @[:@29211.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29213.4]
  assign RetimeWrapper_40_io_in = x460_sum_1_io_result; // @[package.scala 94:16:@29212.4]
  assign x259_div_1_clock = clock; // @[:@29224.4]
  assign x259_div_1_io_a = x254_rdcol_1_io_result; // @[Math.scala 328:17:@29226.4]
  assign x259_div_1_io_flow = io_in_x195_TREADY; // @[Math.scala 330:20:@29228.4]
  assign x260_sum_1_clock = clock; // @[:@29234.4]
  assign x260_sum_1_reset = reset; // @[:@29235.4]
  assign x260_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@29236.4]
  assign x260_sum_1_io_b = x259_div_1_io_result; // @[Math.scala 152:17:@29237.4]
  assign x260_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29238.4]
  assign RetimeWrapper_41_clock = clock; // @[:@29244.4]
  assign RetimeWrapper_41_reset = reset; // @[:@29245.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29247.4]
  assign RetimeWrapper_41_io_in = ~ x256; // @[package.scala 94:16:@29246.4]
  assign RetimeWrapper_42_clock = clock; // @[:@29253.4]
  assign RetimeWrapper_42_reset = reset; // @[:@29254.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29256.4]
  assign RetimeWrapper_42_io_in = x461 ? x503_x460_sum_D1_number : x463_sub_number; // @[package.scala 94:16:@29255.4]
  assign RetimeWrapper_43_clock = clock; // @[:@29265.4]
  assign RetimeWrapper_43_reset = reset; // @[:@29266.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29268.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29267.4]
  assign x263_rdrow_1_clock = clock; // @[:@29288.4]
  assign x263_rdrow_1_reset = reset; // @[:@29289.4]
  assign x263_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@29290.4]
  assign x263_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@29291.4]
  assign x263_rdrow_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@29292.4]
  assign RetimeWrapper_44_clock = clock; // @[:@29314.4]
  assign RetimeWrapper_44_reset = reset; // @[:@29315.4]
  assign RetimeWrapper_44_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29317.4]
  assign RetimeWrapper_44_io_in = $signed(_T_1393) < $signed(32'sh0); // @[package.scala 94:16:@29316.4]
  assign RetimeWrapper_45_clock = clock; // @[:@29323.4]
  assign RetimeWrapper_45_reset = reset; // @[:@29324.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29326.4]
  assign RetimeWrapper_45_io_in = RetimeWrapper_16_io_out; // @[package.scala 94:16:@29325.4]
  assign RetimeWrapper_46_clock = clock; // @[:@29345.4]
  assign RetimeWrapper_46_reset = reset; // @[:@29346.4]
  assign RetimeWrapper_46_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29349.4]
  assign RetimeWrapper_46_io_in = $unsigned(_T_1425); // @[package.scala 94:16:@29348.4]
  assign RetimeWrapper_47_clock = clock; // @[:@29371.4]
  assign RetimeWrapper_47_reset = reset; // @[:@29372.4]
  assign RetimeWrapper_47_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29374.4]
  assign RetimeWrapper_47_io_in = {_T_1437,_T_1438}; // @[package.scala 94:16:@29373.4]
  assign x469_sum_1_clock = clock; // @[:@29392.4]
  assign x469_sum_1_reset = reset; // @[:@29393.4]
  assign x469_sum_1_io_a = _T_1461[31:0]; // @[Math.scala 151:17:@29394.4]
  assign x469_sum_1_io_b = _T_1464[31:0]; // @[Math.scala 152:17:@29395.4]
  assign x469_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29396.4]
  assign RetimeWrapper_48_clock = clock; // @[:@29402.4]
  assign RetimeWrapper_48_reset = reset; // @[:@29403.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29405.4]
  assign RetimeWrapper_48_io_in = x469_sum_1_io_result; // @[package.scala 94:16:@29404.4]
  assign RetimeWrapper_49_clock = clock; // @[:@29411.4]
  assign RetimeWrapper_49_reset = reset; // @[:@29412.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29414.4]
  assign RetimeWrapper_49_io_in = x235_div_1_io_result; // @[package.scala 94:16:@29413.4]
  assign x271_sum_1_clock = clock; // @[:@29420.4]
  assign x271_sum_1_reset = reset; // @[:@29421.4]
  assign x271_sum_1_io_a = RetimeWrapper_48_io_out; // @[Math.scala 151:17:@29422.4]
  assign x271_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@29423.4]
  assign x271_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29424.4]
  assign RetimeWrapper_50_clock = clock; // @[:@29430.4]
  assign RetimeWrapper_50_reset = reset; // @[:@29431.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29433.4]
  assign RetimeWrapper_50_io_in = $unsigned(_T_1429); // @[package.scala 94:16:@29432.4]
  assign RetimeWrapper_51_clock = clock; // @[:@29439.4]
  assign RetimeWrapper_51_reset = reset; // @[:@29440.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29442.4]
  assign RetimeWrapper_51_io_in = x271_sum_1_io_result; // @[package.scala 94:16:@29441.4]
  assign RetimeWrapper_52_clock = clock; // @[:@29448.4]
  assign RetimeWrapper_52_reset = reset; // @[:@29449.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29451.4]
  assign RetimeWrapper_52_io_in = ~ x266; // @[package.scala 94:16:@29450.4]
  assign RetimeWrapper_53_clock = clock; // @[:@29460.4]
  assign RetimeWrapper_53_reset = reset; // @[:@29461.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29463.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29462.4]
  assign RetimeWrapper_54_clock = clock; // @[:@29487.4]
  assign RetimeWrapper_54_reset = reset; // @[:@29488.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29490.4]
  assign RetimeWrapper_54_io_in = x469_sum_1_io_result; // @[package.scala 94:16:@29489.4]
  assign x276_sum_1_clock = clock; // @[:@29498.4]
  assign x276_sum_1_reset = reset; // @[:@29499.4]
  assign x276_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@29500.4]
  assign x276_sum_1_io_b = x250_div_1_io_result; // @[Math.scala 152:17:@29501.4]
  assign x276_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29502.4]
  assign RetimeWrapper_55_clock = clock; // @[:@29508.4]
  assign RetimeWrapper_55_reset = reset; // @[:@29509.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29511.4]
  assign RetimeWrapper_55_io_in = ~ x274; // @[package.scala 94:16:@29510.4]
  assign RetimeWrapper_56_clock = clock; // @[:@29520.4]
  assign RetimeWrapper_56_reset = reset; // @[:@29521.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29523.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29522.4]
  assign x281_sum_1_clock = clock; // @[:@29547.4]
  assign x281_sum_1_reset = reset; // @[:@29548.4]
  assign x281_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@29549.4]
  assign x281_sum_1_io_b = x259_div_1_io_result; // @[Math.scala 152:17:@29550.4]
  assign x281_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29551.4]
  assign RetimeWrapper_57_clock = clock; // @[:@29557.4]
  assign RetimeWrapper_57_reset = reset; // @[:@29558.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29560.4]
  assign RetimeWrapper_57_io_in = ~ x279; // @[package.scala 94:16:@29559.4]
  assign RetimeWrapper_58_clock = clock; // @[:@29569.4]
  assign RetimeWrapper_58_reset = reset; // @[:@29570.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29572.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29571.4]
  assign x284_rdrow_1_clock = clock; // @[:@29592.4]
  assign x284_rdrow_1_reset = reset; // @[:@29593.4]
  assign x284_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@29594.4]
  assign x284_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@29595.4]
  assign x284_rdrow_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@29596.4]
  assign RetimeWrapper_59_clock = clock; // @[:@29618.4]
  assign RetimeWrapper_59_reset = reset; // @[:@29619.4]
  assign RetimeWrapper_59_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29621.4]
  assign RetimeWrapper_59_io_in = $signed(_T_1582) < $signed(32'sh0); // @[package.scala 94:16:@29620.4]
  assign RetimeWrapper_60_clock = clock; // @[:@29640.4]
  assign RetimeWrapper_60_reset = reset; // @[:@29641.4]
  assign RetimeWrapper_60_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29644.4]
  assign RetimeWrapper_60_io_in = $unsigned(_T_1611); // @[package.scala 94:16:@29643.4]
  assign RetimeWrapper_61_clock = clock; // @[:@29666.4]
  assign RetimeWrapper_61_reset = reset; // @[:@29667.4]
  assign RetimeWrapper_61_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@29669.4]
  assign RetimeWrapper_61_io_in = {_T_1623,_T_1624}; // @[package.scala 94:16:@29668.4]
  assign x474_sum_1_clock = clock; // @[:@29687.4]
  assign x474_sum_1_reset = reset; // @[:@29688.4]
  assign x474_sum_1_io_a = _T_1647[31:0]; // @[Math.scala 151:17:@29689.4]
  assign x474_sum_1_io_b = _T_1650[31:0]; // @[Math.scala 152:17:@29690.4]
  assign x474_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29691.4]
  assign RetimeWrapper_62_clock = clock; // @[:@29697.4]
  assign RetimeWrapper_62_reset = reset; // @[:@29698.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29700.4]
  assign RetimeWrapper_62_io_in = x474_sum_1_io_result; // @[package.scala 94:16:@29699.4]
  assign x292_sum_1_clock = clock; // @[:@29706.4]
  assign x292_sum_1_reset = reset; // @[:@29707.4]
  assign x292_sum_1_io_a = RetimeWrapper_62_io_out; // @[Math.scala 151:17:@29708.4]
  assign x292_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@29709.4]
  assign x292_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29710.4]
  assign RetimeWrapper_63_clock = clock; // @[:@29716.4]
  assign RetimeWrapper_63_reset = reset; // @[:@29717.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29719.4]
  assign RetimeWrapper_63_io_in = ~ x287; // @[package.scala 94:16:@29718.4]
  assign RetimeWrapper_64_clock = clock; // @[:@29725.4]
  assign RetimeWrapper_64_reset = reset; // @[:@29726.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29728.4]
  assign RetimeWrapper_64_io_in = x292_sum_1_io_result; // @[package.scala 94:16:@29727.4]
  assign RetimeWrapper_65_clock = clock; // @[:@29734.4]
  assign RetimeWrapper_65_reset = reset; // @[:@29735.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29737.4]
  assign RetimeWrapper_65_io_in = $unsigned(_T_1615); // @[package.scala 94:16:@29736.4]
  assign RetimeWrapper_66_clock = clock; // @[:@29746.4]
  assign RetimeWrapper_66_reset = reset; // @[:@29747.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29749.4]
  assign RetimeWrapper_66_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29748.4]
  assign RetimeWrapper_67_clock = clock; // @[:@29773.4]
  assign RetimeWrapper_67_reset = reset; // @[:@29774.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29776.4]
  assign RetimeWrapper_67_io_in = x474_sum_1_io_result; // @[package.scala 94:16:@29775.4]
  assign x297_sum_1_clock = clock; // @[:@29782.4]
  assign x297_sum_1_reset = reset; // @[:@29783.4]
  assign x297_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@29784.4]
  assign x297_sum_1_io_b = x250_div_1_io_result; // @[Math.scala 152:17:@29785.4]
  assign x297_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29786.4]
  assign RetimeWrapper_68_clock = clock; // @[:@29792.4]
  assign RetimeWrapper_68_reset = reset; // @[:@29793.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29795.4]
  assign RetimeWrapper_68_io_in = ~ x295; // @[package.scala 94:16:@29794.4]
  assign RetimeWrapper_69_clock = clock; // @[:@29804.4]
  assign RetimeWrapper_69_reset = reset; // @[:@29805.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29807.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29806.4]
  assign x302_sum_1_clock = clock; // @[:@29831.4]
  assign x302_sum_1_reset = reset; // @[:@29832.4]
  assign x302_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@29833.4]
  assign x302_sum_1_io_b = x259_div_1_io_result; // @[Math.scala 152:17:@29834.4]
  assign x302_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29835.4]
  assign RetimeWrapper_70_clock = clock; // @[:@29841.4]
  assign RetimeWrapper_70_reset = reset; // @[:@29842.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29844.4]
  assign RetimeWrapper_70_io_in = ~ x300; // @[package.scala 94:16:@29843.4]
  assign RetimeWrapper_71_clock = clock; // @[:@29853.4]
  assign RetimeWrapper_71_reset = reset; // @[:@29854.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29856.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29855.4]
  assign x305_1_clock = clock; // @[:@29876.4]
  assign x305_1_io_a = x227_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@29878.4]
  assign x305_1_io_b = 32'h1; // @[Math.scala 264:17:@29879.4]
  assign x305_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29880.4]
  assign x306_1_clock = clock; // @[:@29888.4]
  assign x306_1_io_a = x227_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@29890.4]
  assign x306_1_io_b = 32'h2; // @[Math.scala 264:17:@29891.4]
  assign x306_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29892.4]
  assign x307_1_clock = clock; // @[:@29900.4]
  assign x307_1_io_a = x227_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@29902.4]
  assign x307_1_io_b = 32'h1; // @[Math.scala 264:17:@29903.4]
  assign x307_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29904.4]
  assign x308_1_clock = clock; // @[:@29912.4]
  assign x308_1_io_a = x227_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@29914.4]
  assign x308_1_io_b = 32'h2; // @[Math.scala 264:17:@29915.4]
  assign x308_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29916.4]
  assign x309_1_clock = clock; // @[:@29924.4]
  assign x309_1_io_a = x227_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@29926.4]
  assign x309_1_io_b = 32'h4; // @[Math.scala 264:17:@29927.4]
  assign x309_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29928.4]
  assign x310_1_clock = clock; // @[:@29938.4]
  assign x310_1_io_a = x227_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@29940.4]
  assign x310_1_io_b = 32'h2; // @[Math.scala 264:17:@29941.4]
  assign x310_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29942.4]
  assign x311_1_clock = clock; // @[:@29950.4]
  assign x311_1_io_a = x227_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@29952.4]
  assign x311_1_io_b = 32'h1; // @[Math.scala 264:17:@29953.4]
  assign x311_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29954.4]
  assign x312_1_clock = clock; // @[:@29962.4]
  assign x312_1_io_a = x227_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@29964.4]
  assign x312_1_io_b = 32'h2; // @[Math.scala 264:17:@29965.4]
  assign x312_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29966.4]
  assign x313_1_clock = clock; // @[:@29974.4]
  assign x313_1_io_a = x227_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@29976.4]
  assign x313_1_io_b = 32'h1; // @[Math.scala 264:17:@29977.4]
  assign x313_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@29978.4]
  assign x314_x13_1_clock = clock; // @[:@29984.4]
  assign x314_x13_1_reset = reset; // @[:@29985.4]
  assign x314_x13_1_io_a = x305_1_io_result; // @[Math.scala 151:17:@29986.4]
  assign x314_x13_1_io_b = x306_1_io_result; // @[Math.scala 152:17:@29987.4]
  assign x314_x13_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29988.4]
  assign x315_x14_1_clock = clock; // @[:@29994.4]
  assign x315_x14_1_reset = reset; // @[:@29995.4]
  assign x315_x14_1_io_a = x307_1_io_result; // @[Math.scala 151:17:@29996.4]
  assign x315_x14_1_io_b = x308_1_io_result; // @[Math.scala 152:17:@29997.4]
  assign x315_x14_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@29998.4]
  assign x316_x13_1_clock = clock; // @[:@30004.4]
  assign x316_x13_1_reset = reset; // @[:@30005.4]
  assign x316_x13_1_io_a = x309_1_io_result; // @[Math.scala 151:17:@30006.4]
  assign x316_x13_1_io_b = x310_1_io_result; // @[Math.scala 152:17:@30007.4]
  assign x316_x13_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@30008.4]
  assign x317_x14_1_clock = clock; // @[:@30014.4]
  assign x317_x14_1_reset = reset; // @[:@30015.4]
  assign x317_x14_1_io_a = x311_1_io_result; // @[Math.scala 151:17:@30016.4]
  assign x317_x14_1_io_b = x312_1_io_result; // @[Math.scala 152:17:@30017.4]
  assign x317_x14_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@30018.4]
  assign x318_x13_1_clock = clock; // @[:@30024.4]
  assign x318_x13_1_reset = reset; // @[:@30025.4]
  assign x318_x13_1_io_a = x314_x13_1_io_result; // @[Math.scala 151:17:@30026.4]
  assign x318_x13_1_io_b = x315_x14_1_io_result; // @[Math.scala 152:17:@30027.4]
  assign x318_x13_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@30028.4]
  assign x319_x14_1_clock = clock; // @[:@30034.4]
  assign x319_x14_1_reset = reset; // @[:@30035.4]
  assign x319_x14_1_io_a = x316_x13_1_io_result; // @[Math.scala 151:17:@30036.4]
  assign x319_x14_1_io_b = x317_x14_1_io_result; // @[Math.scala 152:17:@30037.4]
  assign x319_x14_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@30038.4]
  assign x320_x13_1_clock = clock; // @[:@30044.4]
  assign x320_x13_1_reset = reset; // @[:@30045.4]
  assign x320_x13_1_io_a = x318_x13_1_io_result; // @[Math.scala 151:17:@30046.4]
  assign x320_x13_1_io_b = x319_x14_1_io_result; // @[Math.scala 152:17:@30047.4]
  assign x320_x13_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@30048.4]
  assign RetimeWrapper_72_clock = clock; // @[:@30054.4]
  assign RetimeWrapper_72_reset = reset; // @[:@30055.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30057.4]
  assign RetimeWrapper_72_io_in = x313_1_io_result; // @[package.scala 94:16:@30056.4]
  assign x321_sum_1_clock = clock; // @[:@30063.4]
  assign x321_sum_1_reset = reset; // @[:@30064.4]
  assign x321_sum_1_io_a = x320_x13_1_io_result; // @[Math.scala 151:17:@30065.4]
  assign x321_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@30066.4]
  assign x321_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@30067.4]
  assign x322_1_io_b = x321_sum_1_io_result; // @[Math.scala 721:17:@30075.4]
  assign x323_mul_1_clock = clock; // @[:@30084.4]
  assign x323_mul_1_io_a = x322_1_io_result; // @[Math.scala 263:17:@30086.4]
  assign x323_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@30087.4]
  assign x323_mul_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@30088.4]
  assign x324_1_io_b = x323_mul_1_io_result; // @[Math.scala 721:17:@30096.4]
  assign RetimeWrapper_73_clock = clock; // @[:@30103.4]
  assign RetimeWrapper_73_reset = reset; // @[:@30104.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30106.4]
  assign RetimeWrapper_73_io_in = x227_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@30105.4]
  assign x325_sub_1_clock = clock; // @[:@30112.4]
  assign x325_sub_1_reset = reset; // @[:@30113.4]
  assign x325_sub_1_io_a = RetimeWrapper_73_io_out; // @[Math.scala 192:17:@30114.4]
  assign x325_sub_1_io_b = x324_1_io_result; // @[Math.scala 193:17:@30115.4]
  assign x325_sub_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@30116.4]
  assign RetimeWrapper_74_clock = clock; // @[:@30125.4]
  assign RetimeWrapper_74_reset = reset; // @[:@30126.4]
  assign RetimeWrapper_74_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@30128.4]
  assign RetimeWrapper_74_io_in = 32'hf < x325_sub_number; // @[package.scala 94:16:@30127.4]
  assign x327_sub_1_clock = clock; // @[:@30134.4]
  assign x327_sub_1_reset = reset; // @[:@30135.4]
  assign x327_sub_1_io_a = x324_1_io_result; // @[Math.scala 192:17:@30136.4]
  assign x327_sub_1_io_b = RetimeWrapper_73_io_out; // @[Math.scala 193:17:@30137.4]
  assign x327_sub_1_io_flow = io_in_x195_TREADY; // @[Math.scala 194:20:@30138.4]
  assign RetimeWrapper_75_clock = clock; // @[:@30147.4]
  assign RetimeWrapper_75_reset = reset; // @[:@30148.4]
  assign RetimeWrapper_75_io_flow = io_in_x195_TREADY; // @[package.scala 95:18:@30150.4]
  assign RetimeWrapper_75_io_in = 32'hf < x327_sub_number; // @[package.scala 94:16:@30149.4]
  assign RetimeWrapper_76_clock = clock; // @[:@30159.4]
  assign RetimeWrapper_76_reset = reset; // @[:@30160.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30162.4]
  assign RetimeWrapper_76_io_in = x325_sub_1_io_result; // @[package.scala 94:16:@30161.4]
  assign x331_1_io_b = x329 ? x524_x325_sub_D1_number : 32'h0; // @[Math.scala 721:17:@30175.4]
  assign x332_mul_1_clock = clock; // @[:@30184.4]
  assign x332_mul_1_io_a = x331_1_io_result; // @[Math.scala 263:17:@30186.4]
  assign x332_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@30187.4]
  assign x332_mul_1_io_flow = io_in_x195_TREADY; // @[Math.scala 265:20:@30188.4]
  assign x333_1_io_b = x332_mul_1_io_result; // @[Math.scala 721:17:@30196.4]
  assign RetimeWrapper_77_clock = clock; // @[:@30203.4]
  assign RetimeWrapper_77_reset = reset; // @[:@30204.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30206.4]
  assign RetimeWrapper_77_io_in = x227_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@30205.4]
  assign x334_sum_1_clock = clock; // @[:@30212.4]
  assign x334_sum_1_reset = reset; // @[:@30213.4]
  assign x334_sum_1_io_a = RetimeWrapper_77_io_out; // @[Math.scala 151:17:@30214.4]
  assign x334_sum_1_io_b = x333_1_io_result; // @[Math.scala 152:17:@30215.4]
  assign x334_sum_1_io_flow = io_in_x195_TREADY; // @[Math.scala 153:20:@30216.4]
  assign RetimeWrapper_78_clock = clock; // @[:@30226.4]
  assign RetimeWrapper_78_reset = reset; // @[:@30227.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30229.4]
  assign RetimeWrapper_78_io_in = x334_sum_1_io_result; // @[package.scala 94:16:@30228.4]
  assign RetimeWrapper_79_clock = clock; // @[:@30235.4]
  assign RetimeWrapper_79_reset = reset; // @[:@30236.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30238.4]
  assign RetimeWrapper_79_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@30237.4]
  assign RetimeWrapper_80_clock = clock; // @[:@30244.4]
  assign RetimeWrapper_80_reset = reset; // @[:@30245.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30247.4]
  assign RetimeWrapper_80_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@30246.4]
  assign RetimeWrapper_81_clock = clock; // @[:@30253.4]
  assign RetimeWrapper_81_reset = reset; // @[:@30254.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30256.4]
  assign RetimeWrapper_81_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@30255.4]
endmodule
module x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1( // @[:@30274.2]
  input          clock, // @[:@30275.4]
  input          reset, // @[:@30276.4]
  input          io_in_x194_TVALID, // @[:@30277.4]
  output         io_in_x194_TREADY, // @[:@30277.4]
  input  [255:0] io_in_x194_TDATA, // @[:@30277.4]
  input  [7:0]   io_in_x194_TID, // @[:@30277.4]
  input  [7:0]   io_in_x194_TDEST, // @[:@30277.4]
  output         io_in_x195_TVALID, // @[:@30277.4]
  input          io_in_x195_TREADY, // @[:@30277.4]
  output [255:0] io_in_x195_TDATA, // @[:@30277.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@30277.4]
  input          io_sigsIn_smChildAcks_0, // @[:@30277.4]
  output         io_sigsOut_smDoneIn_0, // @[:@30277.4]
  input          io_rr // @[:@30277.4]
);
  wire  x220_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire  x220_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire  x220_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire  x220_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire [12:0] x220_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire [12:0] x220_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire  x220_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire  x220_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire  x220_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@30311.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30399.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30399.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30399.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30399.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30399.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30441.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30441.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30441.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30441.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30441.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30449.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30449.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30449.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30449.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30449.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TREADY; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire [255:0] x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TDATA; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire [7:0] x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TID; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire [7:0] x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TDEST; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TVALID; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TREADY; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire [255:0] x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TDATA; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire [31:0] x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire [31:0] x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
  wire  _T_240; // @[package.scala 96:25:@30404.4 package.scala 96:25:@30405.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x340_outr_UnitPipe.scala 69:66:@30410.4]
  wire  _T_253; // @[package.scala 96:25:@30446.4 package.scala 96:25:@30447.4]
  wire  _T_259; // @[package.scala 96:25:@30454.4 package.scala 96:25:@30455.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@30457.4]
  wire  x339_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@30458.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@30466.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@30467.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@30479.4]
  x202_ctrchain x220_ctrchain ( // @[SpatialBlocks.scala 37:22:@30311.4]
    .clock(x220_ctrchain_clock),
    .reset(x220_ctrchain_reset),
    .io_input_reset(x220_ctrchain_io_input_reset),
    .io_input_enable(x220_ctrchain_io_input_enable),
    .io_output_counts_1(x220_ctrchain_io_output_counts_1),
    .io_output_counts_0(x220_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x220_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x220_ctrchain_io_output_oobs_1),
    .io_output_done(x220_ctrchain_io_output_done)
  );
  x339_inr_Foreach_SAMPLER_BOX_sm x339_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 32:18:@30371.4]
    .clock(x339_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x339_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x339_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x339_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x339_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x339_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x339_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x339_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x339_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30399.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30441.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30449.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1 x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 602:24:@30483.4]
    .clock(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x194_TREADY(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TREADY),
    .io_in_x194_TDATA(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TDATA),
    .io_in_x194_TID(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TID),
    .io_in_x194_TDEST(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TDEST),
    .io_in_x195_TVALID(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TVALID),
    .io_in_x195_TREADY(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TREADY),
    .io_in_x195_TDATA(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TDATA),
    .io_sigsIn_backpressure(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@30404.4 package.scala 96:25:@30405.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x194_TVALID | x339_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x340_outr_UnitPipe.scala 69:66:@30410.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30446.4 package.scala 96:25:@30447.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@30454.4 package.scala 96:25:@30455.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@30457.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@30458.4]
  assign _T_264 = x339_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@30466.4]
  assign _T_265 = ~ x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@30467.4]
  assign _T_272 = x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@30479.4]
  assign io_in_x194_TREADY = x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TREADY; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 48:23:@30541.4]
  assign io_in_x195_TVALID = x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TVALID; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 49:23:@30551.4]
  assign io_in_x195_TDATA = x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TDATA; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 49:23:@30549.4]
  assign io_sigsOut_smDoneIn_0 = x339_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@30464.4]
  assign x220_ctrchain_clock = clock; // @[:@30312.4]
  assign x220_ctrchain_reset = reset; // @[:@30313.4]
  assign x220_ctrchain_io_input_reset = x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@30482.4]
  assign x220_ctrchain_io_input_enable = _T_272 & x339_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@30434.4 SpatialBlocks.scala 159:42:@30481.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@30372.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@30373.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sm_io_enable = x339_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x339_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@30461.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x340_outr_UnitPipe.scala 67:50:@30407.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@30463.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x195_TREADY | x339_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@30435.4]
  assign x339_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x340_outr_UnitPipe.scala 71:48:@30413.4]
  assign RetimeWrapper_clock = clock; // @[:@30400.4]
  assign RetimeWrapper_reset = reset; // @[:@30401.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30403.4]
  assign RetimeWrapper_io_in = x220_ctrchain_io_output_done; // @[package.scala 94:16:@30402.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30442.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30443.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30445.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@30444.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30450.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30451.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30453.4]
  assign RetimeWrapper_2_io_in = x339_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@30452.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@30484.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@30485.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TDATA = io_in_x194_TDATA; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 48:23:@30540.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TID = io_in_x194_TID; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 48:23:@30536.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x194_TDEST = io_in_x194_TDEST; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 48:23:@30535.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x195_TREADY = io_in_x195_TREADY; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 49:23:@30550.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x195_TREADY | x339_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 607:22:@30568.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 607:22:@30566.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x339_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 607:22:@30564.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x220_ctrchain_io_output_counts_1[12]}},x220_ctrchain_io_output_counts_1}; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 607:22:@30559.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x220_ctrchain_io_output_counts_0[12]}},x220_ctrchain_io_output_counts_0}; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 607:22:@30558.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x220_ctrchain_io_output_oobs_0; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 607:22:@30556.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x220_ctrchain_io_output_oobs_1; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 607:22:@30557.4]
  assign x339_inr_Foreach_SAMPLER_BOX_kernelx339_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x339_inr_Foreach_SAMPLER_BOX.scala 606:18:@30552.4]
endmodule
module x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1( // @[:@30582.2]
  input          clock, // @[:@30583.4]
  input          reset, // @[:@30584.4]
  input          io_in_x194_TVALID, // @[:@30585.4]
  output         io_in_x194_TREADY, // @[:@30585.4]
  input  [255:0] io_in_x194_TDATA, // @[:@30585.4]
  input  [7:0]   io_in_x194_TID, // @[:@30585.4]
  input  [7:0]   io_in_x194_TDEST, // @[:@30585.4]
  output         io_in_x195_TVALID, // @[:@30585.4]
  input          io_in_x195_TREADY, // @[:@30585.4]
  output [255:0] io_in_x195_TDATA, // @[:@30585.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@30585.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@30585.4]
  input          io_sigsIn_smChildAcks_0, // @[:@30585.4]
  input          io_sigsIn_smChildAcks_1, // @[:@30585.4]
  output         io_sigsOut_smDoneIn_0, // @[:@30585.4]
  output         io_sigsOut_smDoneIn_1, // @[:@30585.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@30585.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@30585.4]
  input          io_rr // @[:@30585.4]
);
  wire  x197_fifoinraw_0_clock; // @[m_x197_fifoinraw_0.scala 27:17:@30599.4]
  wire  x197_fifoinraw_0_reset; // @[m_x197_fifoinraw_0.scala 27:17:@30599.4]
  wire  x198_fifoinpacked_0_clock; // @[m_x198_fifoinpacked_0.scala 27:17:@30623.4]
  wire  x198_fifoinpacked_0_reset; // @[m_x198_fifoinpacked_0.scala 27:17:@30623.4]
  wire  x198_fifoinpacked_0_io_wPort_0_en_0; // @[m_x198_fifoinpacked_0.scala 27:17:@30623.4]
  wire  x198_fifoinpacked_0_io_full; // @[m_x198_fifoinpacked_0.scala 27:17:@30623.4]
  wire  x198_fifoinpacked_0_io_active_0_in; // @[m_x198_fifoinpacked_0.scala 27:17:@30623.4]
  wire  x198_fifoinpacked_0_io_active_0_out; // @[m_x198_fifoinpacked_0.scala 27:17:@30623.4]
  wire  x199_fifooutraw_0_clock; // @[m_x199_fifooutraw_0.scala 27:17:@30647.4]
  wire  x199_fifooutraw_0_reset; // @[m_x199_fifooutraw_0.scala 27:17:@30647.4]
  wire  x202_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire  x202_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire  x202_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire  x202_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire [12:0] x202_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire [12:0] x202_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire  x202_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire  x202_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire  x202_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@30671.4]
  wire  x216_inr_Foreach_sm_clock; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_reset; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_enable; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_done; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_doneLatch; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_ctrDone; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_datapathEn; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_ctrInc; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_ctrRst; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_parentAck; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_backpressure; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  x216_inr_Foreach_sm_io_break; // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30759.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30759.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30759.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30759.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30759.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30805.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30805.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30805.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30805.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30805.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30813.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30813.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30813.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30813.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30813.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_clock; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_reset; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_wPort_0_en_0; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_full; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_active_0_in; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_active_0_out; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire [31:0] x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire [31:0] x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_rr; // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
  wire  x340_outr_UnitPipe_sm_clock; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_reset; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_enable; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_done; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_rst; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_ctrDone; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_ctrInc; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_parentAck; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  x340_outr_UnitPipe_sm_io_childAck_0; // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31037.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31037.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31037.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31037.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31037.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@31045.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@31045.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@31045.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@31045.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@31045.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_clock; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_reset; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TVALID; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TREADY; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire [255:0] x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TDATA; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire [7:0] x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TID; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire [7:0] x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TDEST; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TVALID; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TREADY; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire [255:0] x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TDATA; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_rr; // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
  wire  _T_254; // @[package.scala 96:25:@30764.4 package.scala 96:25:@30765.4]
  wire  _T_260; // @[implicits.scala 47:10:@30768.4]
  wire  _T_261; // @[sm_x341_outr_UnitPipe.scala 70:41:@30769.4]
  wire  _T_262; // @[sm_x341_outr_UnitPipe.scala 70:78:@30770.4]
  wire  _T_263; // @[sm_x341_outr_UnitPipe.scala 70:76:@30771.4]
  wire  _T_275; // @[package.scala 96:25:@30810.4 package.scala 96:25:@30811.4]
  wire  _T_281; // @[package.scala 96:25:@30818.4 package.scala 96:25:@30819.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@30821.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@30830.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@30831.4]
  wire  _T_354; // @[package.scala 100:49:@31008.4]
  reg  _T_357; // @[package.scala 48:56:@31009.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@31042.4 package.scala 96:25:@31043.4]
  wire  _T_377; // @[package.scala 96:25:@31050.4 package.scala 96:25:@31051.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@31053.4]
  x197_fifoinraw_0 x197_fifoinraw_0 ( // @[m_x197_fifoinraw_0.scala 27:17:@30599.4]
    .clock(x197_fifoinraw_0_clock),
    .reset(x197_fifoinraw_0_reset)
  );
  x198_fifoinpacked_0 x198_fifoinpacked_0 ( // @[m_x198_fifoinpacked_0.scala 27:17:@30623.4]
    .clock(x198_fifoinpacked_0_clock),
    .reset(x198_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x198_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x198_fifoinpacked_0_io_full),
    .io_active_0_in(x198_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x198_fifoinpacked_0_io_active_0_out)
  );
  x197_fifoinraw_0 x199_fifooutraw_0 ( // @[m_x199_fifooutraw_0.scala 27:17:@30647.4]
    .clock(x199_fifooutraw_0_clock),
    .reset(x199_fifooutraw_0_reset)
  );
  x202_ctrchain x202_ctrchain ( // @[SpatialBlocks.scala 37:22:@30671.4]
    .clock(x202_ctrchain_clock),
    .reset(x202_ctrchain_reset),
    .io_input_reset(x202_ctrchain_io_input_reset),
    .io_input_enable(x202_ctrchain_io_input_enable),
    .io_output_counts_1(x202_ctrchain_io_output_counts_1),
    .io_output_counts_0(x202_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x202_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x202_ctrchain_io_output_oobs_1),
    .io_output_done(x202_ctrchain_io_output_done)
  );
  x216_inr_Foreach_sm x216_inr_Foreach_sm ( // @[sm_x216_inr_Foreach.scala 32:18:@30731.4]
    .clock(x216_inr_Foreach_sm_clock),
    .reset(x216_inr_Foreach_sm_reset),
    .io_enable(x216_inr_Foreach_sm_io_enable),
    .io_done(x216_inr_Foreach_sm_io_done),
    .io_doneLatch(x216_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x216_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x216_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x216_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x216_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x216_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x216_inr_Foreach_sm_io_backpressure),
    .io_break(x216_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30759.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30805.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30813.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x216_inr_Foreach_kernelx216_inr_Foreach_concrete1 x216_inr_Foreach_kernelx216_inr_Foreach_concrete1 ( // @[sm_x216_inr_Foreach.scala 96:24:@30848.4]
    .clock(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_clock),
    .reset(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_reset),
    .io_in_x198_fifoinpacked_0_wPort_0_en_0(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_wPort_0_en_0),
    .io_in_x198_fifoinpacked_0_full(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_full),
    .io_in_x198_fifoinpacked_0_active_0_in(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_active_0_in),
    .io_in_x198_fifoinpacked_0_active_0_out(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x340_outr_UnitPipe_sm ( // @[sm_x340_outr_UnitPipe.scala 32:18:@30980.4]
    .clock(x340_outr_UnitPipe_sm_clock),
    .reset(x340_outr_UnitPipe_sm_reset),
    .io_enable(x340_outr_UnitPipe_sm_io_enable),
    .io_done(x340_outr_UnitPipe_sm_io_done),
    .io_rst(x340_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x340_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x340_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x340_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x340_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x340_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x340_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31037.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@31045.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1 x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1 ( // @[sm_x340_outr_UnitPipe.scala 76:24:@31075.4]
    .clock(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_clock),
    .reset(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_reset),
    .io_in_x194_TVALID(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TVALID),
    .io_in_x194_TREADY(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TREADY),
    .io_in_x194_TDATA(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TDATA),
    .io_in_x194_TID(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TID),
    .io_in_x194_TDEST(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TDEST),
    .io_in_x195_TVALID(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TVALID),
    .io_in_x195_TREADY(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TREADY),
    .io_in_x195_TDATA(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TDATA),
    .io_sigsIn_smEnableOuts_0(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@30764.4 package.scala 96:25:@30765.4]
  assign _T_260 = x198_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@30768.4]
  assign _T_261 = ~ _T_260; // @[sm_x341_outr_UnitPipe.scala 70:41:@30769.4]
  assign _T_262 = ~ x198_fifoinpacked_0_io_active_0_out; // @[sm_x341_outr_UnitPipe.scala 70:78:@30770.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x341_outr_UnitPipe.scala 70:76:@30771.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30810.4 package.scala 96:25:@30811.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@30818.4 package.scala 96:25:@30819.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@30821.4]
  assign _T_286 = x216_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@30830.4]
  assign _T_287 = ~ x216_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@30831.4]
  assign _T_354 = x340_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@31008.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@31042.4 package.scala 96:25:@31043.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@31050.4 package.scala 96:25:@31051.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@31053.4]
  assign io_in_x194_TREADY = x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TREADY; // @[sm_x340_outr_UnitPipe.scala 48:23:@31131.4]
  assign io_in_x195_TVALID = x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TVALID; // @[sm_x340_outr_UnitPipe.scala 49:23:@31141.4]
  assign io_in_x195_TDATA = x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TDATA; // @[sm_x340_outr_UnitPipe.scala 49:23:@31139.4]
  assign io_sigsOut_smDoneIn_0 = x216_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@30828.4]
  assign io_sigsOut_smDoneIn_1 = x340_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@31060.4]
  assign io_sigsOut_smCtrCopyDone_0 = x216_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@30847.4]
  assign io_sigsOut_smCtrCopyDone_1 = x340_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@31074.4]
  assign x197_fifoinraw_0_clock = clock; // @[:@30600.4]
  assign x197_fifoinraw_0_reset = reset; // @[:@30601.4]
  assign x198_fifoinpacked_0_clock = clock; // @[:@30624.4]
  assign x198_fifoinpacked_0_reset = reset; // @[:@30625.4]
  assign x198_fifoinpacked_0_io_wPort_0_en_0 = x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@30908.4]
  assign x198_fifoinpacked_0_io_active_0_in = x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@30907.4]
  assign x199_fifooutraw_0_clock = clock; // @[:@30648.4]
  assign x199_fifooutraw_0_reset = reset; // @[:@30649.4]
  assign x202_ctrchain_clock = clock; // @[:@30672.4]
  assign x202_ctrchain_reset = reset; // @[:@30673.4]
  assign x202_ctrchain_io_input_reset = x216_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@30846.4]
  assign x202_ctrchain_io_input_enable = x216_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@30798.4 SpatialBlocks.scala 159:42:@30845.4]
  assign x216_inr_Foreach_sm_clock = clock; // @[:@30732.4]
  assign x216_inr_Foreach_sm_reset = reset; // @[:@30733.4]
  assign x216_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@30825.4]
  assign x216_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x341_outr_UnitPipe.scala 69:38:@30767.4]
  assign x216_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@30827.4]
  assign x216_inr_Foreach_sm_io_backpressure = _T_263 | x216_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@30799.4]
  assign x216_inr_Foreach_sm_io_break = 1'h0; // @[sm_x341_outr_UnitPipe.scala 73:36:@30777.4]
  assign RetimeWrapper_clock = clock; // @[:@30760.4]
  assign RetimeWrapper_reset = reset; // @[:@30761.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30763.4]
  assign RetimeWrapper_io_in = x202_ctrchain_io_output_done; // @[package.scala 94:16:@30762.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30806.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30807.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30809.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@30808.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30814.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30815.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30817.4]
  assign RetimeWrapper_2_io_in = x216_inr_Foreach_sm_io_done; // @[package.scala 94:16:@30816.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_clock = clock; // @[:@30849.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_reset = reset; // @[:@30850.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_full = x198_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@30902.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_in_x198_fifoinpacked_0_active_0_out = x198_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@30901.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x216_inr_Foreach_sm_io_doneLatch; // @[sm_x216_inr_Foreach.scala 101:22:@30931.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x216_inr_Foreach.scala 101:22:@30929.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_break = x216_inr_Foreach_sm_io_break; // @[sm_x216_inr_Foreach.scala 101:22:@30927.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x202_ctrchain_io_output_counts_1[12]}},x202_ctrchain_io_output_counts_1}; // @[sm_x216_inr_Foreach.scala 101:22:@30922.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x202_ctrchain_io_output_counts_0[12]}},x202_ctrchain_io_output_counts_0}; // @[sm_x216_inr_Foreach.scala 101:22:@30921.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x202_ctrchain_io_output_oobs_0; // @[sm_x216_inr_Foreach.scala 101:22:@30919.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x202_ctrchain_io_output_oobs_1; // @[sm_x216_inr_Foreach.scala 101:22:@30920.4]
  assign x216_inr_Foreach_kernelx216_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x216_inr_Foreach.scala 100:18:@30915.4]
  assign x340_outr_UnitPipe_sm_clock = clock; // @[:@30981.4]
  assign x340_outr_UnitPipe_sm_reset = reset; // @[:@30982.4]
  assign x340_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@31057.4]
  assign x340_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@31032.4]
  assign x340_outr_UnitPipe_sm_io_ctrDone = x340_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x341_outr_UnitPipe.scala 78:40:@31012.4]
  assign x340_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@31059.4]
  assign x340_outr_UnitPipe_sm_io_doneIn_0 = x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@31029.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31038.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31039.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31041.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@31040.4]
  assign RetimeWrapper_4_clock = clock; // @[:@31046.4]
  assign RetimeWrapper_4_reset = reset; // @[:@31047.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@31049.4]
  assign RetimeWrapper_4_io_in = x340_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@31048.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_clock = clock; // @[:@31076.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_reset = reset; // @[:@31077.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TVALID = io_in_x194_TVALID; // @[sm_x340_outr_UnitPipe.scala 48:23:@31132.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TDATA = io_in_x194_TDATA; // @[sm_x340_outr_UnitPipe.scala 48:23:@31130.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TID = io_in_x194_TID; // @[sm_x340_outr_UnitPipe.scala 48:23:@31126.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x194_TDEST = io_in_x194_TDEST; // @[sm_x340_outr_UnitPipe.scala 48:23:@31125.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_in_x195_TREADY = io_in_x195_TREADY; // @[sm_x340_outr_UnitPipe.scala 49:23:@31140.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x340_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x340_outr_UnitPipe.scala 81:22:@31150.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x340_outr_UnitPipe_sm_io_childAck_0; // @[sm_x340_outr_UnitPipe.scala 81:22:@31148.4]
  assign x340_outr_UnitPipe_kernelx340_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x340_outr_UnitPipe.scala 80:18:@31142.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x363_outr_UnitPipe_sm( // @[:@31639.2]
  input   clock, // @[:@31640.4]
  input   reset, // @[:@31641.4]
  input   io_enable, // @[:@31642.4]
  output  io_done, // @[:@31642.4]
  input   io_parentAck, // @[:@31642.4]
  input   io_doneIn_0, // @[:@31642.4]
  input   io_doneIn_1, // @[:@31642.4]
  input   io_doneIn_2, // @[:@31642.4]
  output  io_enableOut_0, // @[:@31642.4]
  output  io_enableOut_1, // @[:@31642.4]
  output  io_enableOut_2, // @[:@31642.4]
  output  io_childAck_0, // @[:@31642.4]
  output  io_childAck_1, // @[:@31642.4]
  output  io_childAck_2, // @[:@31642.4]
  input   io_ctrCopyDone_0, // @[:@31642.4]
  input   io_ctrCopyDone_1, // @[:@31642.4]
  input   io_ctrCopyDone_2 // @[:@31642.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@31645.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@31645.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@31645.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@31645.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@31645.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@31645.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@31648.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@31648.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@31648.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@31648.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@31648.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@31648.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@31651.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@31651.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@31651.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@31651.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@31651.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@31651.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@31654.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@31654.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@31654.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@31654.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@31654.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@31654.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@31657.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@31657.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@31657.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@31657.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@31657.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@31657.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@31660.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@31660.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@31660.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@31660.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@31660.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@31660.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@31701.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@31701.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@31701.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@31701.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@31701.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@31701.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@31704.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@31704.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@31704.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@31704.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@31704.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@31704.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@31707.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@31707.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@31707.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@31707.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@31707.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@31707.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31758.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31758.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31758.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31758.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31758.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31772.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31772.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31772.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31772.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31772.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31790.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31790.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31790.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31790.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31790.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31827.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31827.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31827.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31827.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31827.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@31841.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@31841.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@31841.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@31841.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@31841.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@31859.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@31859.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@31859.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@31859.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@31859.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@31896.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@31896.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@31896.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@31896.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@31896.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@31910.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@31910.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@31910.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@31910.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@31910.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@31985.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@31985.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@31985.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@31985.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@31985.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@32002.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@32002.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@32002.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@32002.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@32002.4]
  wire  _T_77; // @[Controllers.scala 80:47:@31663.4]
  wire  allDone; // @[Controllers.scala 80:47:@31664.4]
  wire  _T_151; // @[Controllers.scala 165:35:@31742.4]
  wire  _T_153; // @[Controllers.scala 165:60:@31743.4]
  wire  _T_154; // @[Controllers.scala 165:58:@31744.4]
  wire  _T_156; // @[Controllers.scala 165:76:@31745.4]
  wire  _T_157; // @[Controllers.scala 165:74:@31746.4]
  wire  _T_161; // @[Controllers.scala 165:109:@31749.4]
  wire  _T_164; // @[Controllers.scala 165:141:@31751.4]
  wire  _T_172; // @[package.scala 96:25:@31763.4 package.scala 96:25:@31764.4]
  wire  _T_176; // @[Controllers.scala 167:54:@31766.4]
  wire  _T_177; // @[Controllers.scala 167:52:@31767.4]
  wire  _T_184; // @[package.scala 96:25:@31777.4 package.scala 96:25:@31778.4]
  wire  _T_202; // @[package.scala 96:25:@31795.4 package.scala 96:25:@31796.4]
  wire  _T_206; // @[Controllers.scala 169:67:@31798.4]
  wire  _T_207; // @[Controllers.scala 169:86:@31799.4]
  wire  _T_219; // @[Controllers.scala 165:35:@31811.4]
  wire  _T_221; // @[Controllers.scala 165:60:@31812.4]
  wire  _T_222; // @[Controllers.scala 165:58:@31813.4]
  wire  _T_224; // @[Controllers.scala 165:76:@31814.4]
  wire  _T_225; // @[Controllers.scala 165:74:@31815.4]
  wire  _T_229; // @[Controllers.scala 165:109:@31818.4]
  wire  _T_232; // @[Controllers.scala 165:141:@31820.4]
  wire  _T_240; // @[package.scala 96:25:@31832.4 package.scala 96:25:@31833.4]
  wire  _T_244; // @[Controllers.scala 167:54:@31835.4]
  wire  _T_245; // @[Controllers.scala 167:52:@31836.4]
  wire  _T_252; // @[package.scala 96:25:@31846.4 package.scala 96:25:@31847.4]
  wire  _T_270; // @[package.scala 96:25:@31864.4 package.scala 96:25:@31865.4]
  wire  _T_274; // @[Controllers.scala 169:67:@31867.4]
  wire  _T_275; // @[Controllers.scala 169:86:@31868.4]
  wire  _T_287; // @[Controllers.scala 165:35:@31880.4]
  wire  _T_289; // @[Controllers.scala 165:60:@31881.4]
  wire  _T_290; // @[Controllers.scala 165:58:@31882.4]
  wire  _T_292; // @[Controllers.scala 165:76:@31883.4]
  wire  _T_293; // @[Controllers.scala 165:74:@31884.4]
  wire  _T_297; // @[Controllers.scala 165:109:@31887.4]
  wire  _T_300; // @[Controllers.scala 165:141:@31889.4]
  wire  _T_308; // @[package.scala 96:25:@31901.4 package.scala 96:25:@31902.4]
  wire  _T_312; // @[Controllers.scala 167:54:@31904.4]
  wire  _T_313; // @[Controllers.scala 167:52:@31905.4]
  wire  _T_320; // @[package.scala 96:25:@31915.4 package.scala 96:25:@31916.4]
  wire  _T_338; // @[package.scala 96:25:@31933.4 package.scala 96:25:@31934.4]
  wire  _T_342; // @[Controllers.scala 169:67:@31936.4]
  wire  _T_343; // @[Controllers.scala 169:86:@31937.4]
  wire  _T_358; // @[Controllers.scala 213:68:@31955.4]
  wire  _T_360; // @[Controllers.scala 213:90:@31957.4]
  wire  _T_362; // @[Controllers.scala 213:132:@31959.4]
  wire  _T_366; // @[Controllers.scala 213:68:@31964.4]
  wire  _T_368; // @[Controllers.scala 213:90:@31966.4]
  wire  _T_374; // @[Controllers.scala 213:68:@31972.4]
  wire  _T_376; // @[Controllers.scala 213:90:@31974.4]
  wire  _T_383; // @[package.scala 100:49:@31980.4]
  reg  _T_386; // @[package.scala 48:56:@31981.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@31983.4]
  reg  _T_400; // @[package.scala 48:56:@31999.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@31645.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@31648.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@31651.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@31654.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@31657.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@31660.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@31701.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@31704.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@31707.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31758.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31772.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31790.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31827.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@31841.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@31859.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@31896.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@31910.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@31928.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@31985.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@32002.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@31663.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@31664.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@31742.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@31743.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@31744.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@31745.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@31746.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@31749.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@31751.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@31763.4 package.scala 96:25:@31764.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@31766.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@31767.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31777.4 package.scala 96:25:@31778.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@31795.4 package.scala 96:25:@31796.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@31798.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@31799.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@31811.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@31812.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@31813.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@31814.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@31815.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@31818.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@31820.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@31832.4 package.scala 96:25:@31833.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@31835.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@31836.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@31846.4 package.scala 96:25:@31847.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@31864.4 package.scala 96:25:@31865.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@31867.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@31868.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@31880.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@31881.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@31882.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@31883.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@31884.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@31887.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@31889.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@31901.4 package.scala 96:25:@31902.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@31904.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@31905.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@31915.4 package.scala 96:25:@31916.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@31933.4 package.scala 96:25:@31934.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@31936.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@31937.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@31955.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@31957.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@31959.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@31964.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@31966.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@31972.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@31974.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@31980.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@31983.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@32009.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@31963.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@31971.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@31979.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@31950.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@31952.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@31954.4]
  assign active_0_clock = clock; // @[:@31646.4]
  assign active_0_reset = reset; // @[:@31647.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@31753.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@31757.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@31667.4]
  assign active_1_clock = clock; // @[:@31649.4]
  assign active_1_reset = reset; // @[:@31650.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@31822.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@31826.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@31668.4]
  assign active_2_clock = clock; // @[:@31652.4]
  assign active_2_reset = reset; // @[:@31653.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@31891.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@31895.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@31669.4]
  assign done_0_clock = clock; // @[:@31655.4]
  assign done_0_reset = reset; // @[:@31656.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@31803.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@31681.4 Controllers.scala 170:32:@31810.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@31670.4]
  assign done_1_clock = clock; // @[:@31658.4]
  assign done_1_reset = reset; // @[:@31659.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@31872.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@31690.4 Controllers.scala 170:32:@31879.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@31671.4]
  assign done_2_clock = clock; // @[:@31661.4]
  assign done_2_reset = reset; // @[:@31662.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@31941.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@31699.4 Controllers.scala 170:32:@31948.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@31672.4]
  assign iterDone_0_clock = clock; // @[:@31702.4]
  assign iterDone_0_reset = reset; // @[:@31703.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@31771.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@31721.4 Controllers.scala 168:36:@31787.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@31710.4]
  assign iterDone_1_clock = clock; // @[:@31705.4]
  assign iterDone_1_reset = reset; // @[:@31706.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@31840.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@31730.4 Controllers.scala 168:36:@31856.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@31711.4]
  assign iterDone_2_clock = clock; // @[:@31708.4]
  assign iterDone_2_reset = reset; // @[:@31709.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@31909.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@31739.4 Controllers.scala 168:36:@31925.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@31712.4]
  assign RetimeWrapper_clock = clock; // @[:@31759.4]
  assign RetimeWrapper_reset = reset; // @[:@31760.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31762.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@31761.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31773.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31774.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31776.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@31775.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31791.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31792.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31794.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@31793.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31828.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31829.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31831.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@31830.4]
  assign RetimeWrapper_4_clock = clock; // @[:@31842.4]
  assign RetimeWrapper_4_reset = reset; // @[:@31843.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@31845.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@31844.4]
  assign RetimeWrapper_5_clock = clock; // @[:@31860.4]
  assign RetimeWrapper_5_reset = reset; // @[:@31861.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@31863.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@31862.4]
  assign RetimeWrapper_6_clock = clock; // @[:@31897.4]
  assign RetimeWrapper_6_reset = reset; // @[:@31898.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@31900.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@31899.4]
  assign RetimeWrapper_7_clock = clock; // @[:@31911.4]
  assign RetimeWrapper_7_reset = reset; // @[:@31912.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@31914.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@31913.4]
  assign RetimeWrapper_8_clock = clock; // @[:@31929.4]
  assign RetimeWrapper_8_reset = reset; // @[:@31930.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@31932.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@31931.4]
  assign RetimeWrapper_9_clock = clock; // @[:@31986.4]
  assign RetimeWrapper_9_reset = reset; // @[:@31987.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@31989.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@31988.4]
  assign RetimeWrapper_10_clock = clock; // @[:@32003.4]
  assign RetimeWrapper_10_reset = reset; // @[:@32004.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@32006.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@32005.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x349_inr_UnitPipe_sm( // @[:@32182.2]
  input   clock, // @[:@32183.4]
  input   reset, // @[:@32184.4]
  input   io_enable, // @[:@32185.4]
  output  io_done, // @[:@32185.4]
  output  io_doneLatch, // @[:@32185.4]
  input   io_ctrDone, // @[:@32185.4]
  output  io_datapathEn, // @[:@32185.4]
  output  io_ctrInc, // @[:@32185.4]
  input   io_parentAck, // @[:@32185.4]
  input   io_backpressure // @[:@32185.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@32187.4]
  wire  active_reset; // @[Controllers.scala 261:22:@32187.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@32187.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@32187.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@32187.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@32187.4]
  wire  done_clock; // @[Controllers.scala 262:20:@32190.4]
  wire  done_reset; // @[Controllers.scala 262:20:@32190.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@32190.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@32190.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@32190.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@32190.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32244.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32244.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32244.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32244.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32244.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32252.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32252.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32252.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32252.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32252.4]
  wire  _T_80; // @[Controllers.scala 264:48:@32195.4]
  wire  _T_81; // @[Controllers.scala 264:46:@32196.4]
  wire  _T_82; // @[Controllers.scala 264:62:@32197.4]
  wire  _T_83; // @[Controllers.scala 264:60:@32198.4]
  wire  _T_100; // @[package.scala 100:49:@32215.4]
  reg  _T_103; // @[package.scala 48:56:@32216.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@32224.4]
  wire  _T_116; // @[Controllers.scala 283:41:@32232.4]
  wire  _T_117; // @[Controllers.scala 283:59:@32233.4]
  wire  _T_119; // @[Controllers.scala 284:37:@32236.4]
  reg  _T_125; // @[package.scala 48:56:@32240.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@32262.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@32265.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@32267.4]
  wire  _T_152; // @[Controllers.scala 292:61:@32268.4]
  wire  _T_153; // @[Controllers.scala 292:24:@32269.4]
  SRFF active ( // @[Controllers.scala 261:22:@32187.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@32190.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32244.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32252.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@32195.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@32196.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@32197.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@32198.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@32215.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@32224.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@32232.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@32233.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@32236.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@32267.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@32268.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@32269.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@32243.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@32271.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@32235.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@32238.4]
  assign active_clock = clock; // @[:@32188.4]
  assign active_reset = reset; // @[:@32189.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@32200.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@32204.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@32205.4]
  assign done_clock = clock; // @[:@32191.4]
  assign done_reset = reset; // @[:@32192.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@32220.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@32213.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@32214.4]
  assign RetimeWrapper_clock = clock; // @[:@32245.4]
  assign RetimeWrapper_reset = reset; // @[:@32246.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32248.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@32247.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32253.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32254.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32256.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@32255.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1( // @[:@32346.2]
  input  [63:0] io_in_x192_outdram_number, // @[:@32349.4]
  output        io_in_x342_valid, // @[:@32349.4]
  output [63:0] io_in_x342_bits_addr, // @[:@32349.4]
  output [31:0] io_in_x342_bits_size, // @[:@32349.4]
  input         io_sigsIn_backpressure, // @[:@32349.4]
  input         io_sigsIn_datapathEn, // @[:@32349.4]
  input         io_rr // @[:@32349.4]
);
  wire [96:0] x346_tuple; // @[Cat.scala 30:58:@32363.4]
  wire  _T_135; // @[implicits.scala 55:10:@32366.4]
  assign x346_tuple = {33'h7e9000,io_in_x192_outdram_number}; // @[Cat.scala 30:58:@32363.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@32366.4]
  assign io_in_x342_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x349_inr_UnitPipe.scala 65:18:@32369.4]
  assign io_in_x342_bits_addr = x346_tuple[63:0]; // @[sm_x349_inr_UnitPipe.scala 66:22:@32371.4]
  assign io_in_x342_bits_size = x346_tuple[95:64]; // @[sm_x349_inr_UnitPipe.scala 67:22:@32373.4]
endmodule
module FF_13( // @[:@32375.2]
  input         clock, // @[:@32376.4]
  input         reset, // @[:@32377.4]
  output [22:0] io_rPort_0_output_0, // @[:@32378.4]
  input  [22:0] io_wPort_0_data_0, // @[:@32378.4]
  input         io_wPort_0_reset, // @[:@32378.4]
  input         io_wPort_0_en_0 // @[:@32378.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@32393.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@32395.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@32396.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@32395.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@32396.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@32398.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@32413.2]
  input         clock, // @[:@32414.4]
  input         reset, // @[:@32415.4]
  input         io_input_reset, // @[:@32416.4]
  input         io_input_enable, // @[:@32416.4]
  output [22:0] io_output_count_0, // @[:@32416.4]
  output        io_output_oobs_0, // @[:@32416.4]
  output        io_output_done // @[:@32416.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@32429.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@32429.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@32429.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@32429.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@32429.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@32429.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@32445.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@32445.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@32445.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@32445.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@32445.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@32445.4]
  wire  _T_36; // @[Counter.scala 264:45:@32448.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@32473.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@32474.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@32475.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@32476.4]
  wire  _T_57; // @[Counter.scala 293:18:@32478.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@32486.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@32489.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@32490.4]
  wire  _T_75; // @[Counter.scala 322:102:@32494.4]
  wire  _T_77; // @[Counter.scala 322:130:@32495.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@32429.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@32445.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@32448.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@32473.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@32474.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@32475.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@32476.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@32478.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@32486.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@32489.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@32490.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@32494.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@32495.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@32493.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@32497.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@32499.4]
  assign bases_0_clock = clock; // @[:@32430.4]
  assign bases_0_reset = reset; // @[:@32431.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@32492.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@32471.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@32472.4]
  assign SRFF_clock = clock; // @[:@32446.4]
  assign SRFF_reset = reset; // @[:@32447.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@32450.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@32452.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@32453.4]
endmodule
module x351_ctrchain( // @[:@32504.2]
  input         clock, // @[:@32505.4]
  input         reset, // @[:@32506.4]
  input         io_input_reset, // @[:@32507.4]
  input         io_input_enable, // @[:@32507.4]
  output [22:0] io_output_counts_0, // @[:@32507.4]
  output        io_output_oobs_0, // @[:@32507.4]
  output        io_output_done // @[:@32507.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@32509.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@32509.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@32509.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@32509.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@32509.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@32509.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@32509.4]
  reg  wasDone; // @[Counter.scala 542:24:@32518.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@32524.4]
  wire  _T_47; // @[Counter.scala 546:80:@32525.4]
  reg  doneLatch; // @[Counter.scala 550:26:@32530.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@32531.4]
  wire  _T_55; // @[Counter.scala 551:19:@32532.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@32509.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@32524.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@32525.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@32531.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@32532.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@32534.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@32536.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@32527.4]
  assign ctrs_0_clock = clock; // @[:@32510.4]
  assign ctrs_0_reset = reset; // @[:@32511.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@32515.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@32516.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x358_inr_Foreach_sm( // @[:@32724.2]
  input   clock, // @[:@32725.4]
  input   reset, // @[:@32726.4]
  input   io_enable, // @[:@32727.4]
  output  io_done, // @[:@32727.4]
  output  io_doneLatch, // @[:@32727.4]
  input   io_ctrDone, // @[:@32727.4]
  output  io_datapathEn, // @[:@32727.4]
  output  io_ctrInc, // @[:@32727.4]
  output  io_ctrRst, // @[:@32727.4]
  input   io_parentAck, // @[:@32727.4]
  input   io_backpressure, // @[:@32727.4]
  input   io_break // @[:@32727.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@32729.4]
  wire  active_reset; // @[Controllers.scala 261:22:@32729.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@32729.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@32729.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@32729.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@32729.4]
  wire  done_clock; // @[Controllers.scala 262:20:@32732.4]
  wire  done_reset; // @[Controllers.scala 262:20:@32732.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@32732.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@32732.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@32732.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@32732.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32766.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32766.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32766.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32766.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32766.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32788.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32788.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32788.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32788.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32788.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32800.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32800.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32800.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32800.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32800.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32808.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32808.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32808.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32808.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32808.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@32824.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@32824.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@32824.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@32824.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@32824.4]
  wire  _T_80; // @[Controllers.scala 264:48:@32737.4]
  wire  _T_81; // @[Controllers.scala 264:46:@32738.4]
  wire  _T_82; // @[Controllers.scala 264:62:@32739.4]
  wire  _T_83; // @[Controllers.scala 264:60:@32740.4]
  wire  _T_100; // @[package.scala 100:49:@32757.4]
  reg  _T_103; // @[package.scala 48:56:@32758.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@32771.4 package.scala 96:25:@32772.4]
  wire  _T_110; // @[package.scala 100:49:@32773.4]
  reg  _T_113; // @[package.scala 48:56:@32774.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@32776.4]
  wire  _T_118; // @[Controllers.scala 283:41:@32781.4]
  wire  _T_119; // @[Controllers.scala 283:59:@32782.4]
  wire  _T_121; // @[Controllers.scala 284:37:@32785.4]
  wire  _T_124; // @[package.scala 96:25:@32793.4 package.scala 96:25:@32794.4]
  wire  _T_126; // @[package.scala 100:49:@32795.4]
  reg  _T_129; // @[package.scala 48:56:@32796.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@32818.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@32820.4]
  reg  _T_153; // @[package.scala 48:56:@32821.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@32829.4 package.scala 96:25:@32830.4]
  wire  _T_158; // @[Controllers.scala 292:61:@32831.4]
  wire  _T_159; // @[Controllers.scala 292:24:@32832.4]
  SRFF active ( // @[Controllers.scala 261:22:@32729.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@32732.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@32766.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@32788.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32800.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32808.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@32824.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@32737.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@32738.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@32739.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@32740.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@32757.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@32771.4 package.scala 96:25:@32772.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@32773.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@32776.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@32781.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@32782.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@32785.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32793.4 package.scala 96:25:@32794.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@32795.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@32820.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@32829.4 package.scala 96:25:@32830.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@32831.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@32832.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@32799.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@32834.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@32784.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@32787.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@32779.4]
  assign active_clock = clock; // @[:@32730.4]
  assign active_reset = reset; // @[:@32731.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@32742.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@32746.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@32747.4]
  assign done_clock = clock; // @[:@32733.4]
  assign done_reset = reset; // @[:@32734.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@32762.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@32755.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@32756.4]
  assign RetimeWrapper_clock = clock; // @[:@32767.4]
  assign RetimeWrapper_reset = reset; // @[:@32768.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@32770.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@32769.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32789.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32790.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@32792.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@32791.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32801.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32802.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32804.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@32803.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32809.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32810.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32812.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@32811.4]
  assign RetimeWrapper_4_clock = clock; // @[:@32825.4]
  assign RetimeWrapper_4_reset = reset; // @[:@32826.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@32828.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@32827.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x358_inr_Foreach_kernelx358_inr_Foreach_concrete1( // @[:@33041.2]
  input         clock, // @[:@33042.4]
  input         reset, // @[:@33043.4]
  output [20:0] io_in_x196_outbuf_0_rPort_0_ofs_0, // @[:@33044.4]
  output        io_in_x196_outbuf_0_rPort_0_en_0, // @[:@33044.4]
  output        io_in_x196_outbuf_0_rPort_0_backpressure, // @[:@33044.4]
  input  [31:0] io_in_x196_outbuf_0_rPort_0_output_0, // @[:@33044.4]
  output        io_in_x343_valid, // @[:@33044.4]
  output [31:0] io_in_x343_bits_wdata_0, // @[:@33044.4]
  output        io_in_x343_bits_wstrb, // @[:@33044.4]
  input         io_sigsIn_backpressure, // @[:@33044.4]
  input         io_sigsIn_datapathEn, // @[:@33044.4]
  input         io_sigsIn_break, // @[:@33044.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@33044.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@33044.4]
  input         io_rr // @[:@33044.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@33071.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@33071.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33100.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33100.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33100.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33100.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33100.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33109.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33109.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33109.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33109.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33109.4]
  wire  b353; // @[sm_x358_inr_Foreach.scala 62:18:@33079.4]
  wire  _T_274; // @[sm_x358_inr_Foreach.scala 67:129:@33083.4]
  wire  _T_278; // @[implicits.scala 55:10:@33086.4]
  wire  _T_279; // @[sm_x358_inr_Foreach.scala 67:146:@33087.4]
  wire [32:0] x356_tuple; // @[Cat.scala 30:58:@33097.4]
  wire  _T_290; // @[package.scala 96:25:@33114.4 package.scala 96:25:@33115.4]
  wire  _T_292; // @[implicits.scala 55:10:@33116.4]
  wire  x528_b353_D2; // @[package.scala 96:25:@33105.4 package.scala 96:25:@33106.4]
  wire  _T_293; // @[sm_x358_inr_Foreach.scala 74:112:@33117.4]
  wire [31:0] b352_number; // @[Math.scala 723:22:@33076.4 Math.scala 724:14:@33077.4]
  _ _ ( // @[Math.scala 720:24:@33071.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@33100.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@33109.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b353 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x358_inr_Foreach.scala 62:18:@33079.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x358_inr_Foreach.scala 67:129:@33083.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@33086.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x358_inr_Foreach.scala 67:146:@33087.4]
  assign x356_tuple = {1'h1,io_in_x196_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@33097.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33114.4 package.scala 96:25:@33115.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@33116.4]
  assign x528_b353_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@33105.4 package.scala 96:25:@33106.4]
  assign _T_293 = _T_292 & x528_b353_D2; // @[sm_x358_inr_Foreach.scala 74:112:@33117.4]
  assign b352_number = __io_result; // @[Math.scala 723:22:@33076.4 Math.scala 724:14:@33077.4]
  assign io_in_x196_outbuf_0_rPort_0_ofs_0 = b352_number[20:0]; // @[MemInterfaceType.scala 107:54:@33090.4]
  assign io_in_x196_outbuf_0_rPort_0_en_0 = _T_279 & b353; // @[MemInterfaceType.scala 110:79:@33092.4]
  assign io_in_x196_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33091.4]
  assign io_in_x343_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x358_inr_Foreach.scala 74:18:@33119.4]
  assign io_in_x343_bits_wdata_0 = x356_tuple[31:0]; // @[sm_x358_inr_Foreach.scala 75:26:@33121.4]
  assign io_in_x343_bits_wstrb = x356_tuple[32]; // @[sm_x358_inr_Foreach.scala 76:23:@33123.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@33074.4]
  assign RetimeWrapper_clock = clock; // @[:@33101.4]
  assign RetimeWrapper_reset = reset; // @[:@33102.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33104.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33103.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33110.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33111.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33113.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33112.4]
endmodule
module x362_inr_UnitPipe_sm( // @[:@33279.2]
  input   clock, // @[:@33280.4]
  input   reset, // @[:@33281.4]
  input   io_enable, // @[:@33282.4]
  output  io_done, // @[:@33282.4]
  output  io_doneLatch, // @[:@33282.4]
  input   io_ctrDone, // @[:@33282.4]
  output  io_datapathEn, // @[:@33282.4]
  output  io_ctrInc, // @[:@33282.4]
  input   io_parentAck // @[:@33282.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@33284.4]
  wire  active_reset; // @[Controllers.scala 261:22:@33284.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@33284.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@33284.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@33284.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@33284.4]
  wire  done_clock; // @[Controllers.scala 262:20:@33287.4]
  wire  done_reset; // @[Controllers.scala 262:20:@33287.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@33287.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@33287.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@33287.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@33287.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33321.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33321.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33321.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33321.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33321.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33343.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@33355.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@33355.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@33355.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@33355.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@33355.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@33363.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@33363.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@33363.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@33363.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@33363.4]
  wire  _T_80; // @[Controllers.scala 264:48:@33292.4]
  wire  _T_81; // @[Controllers.scala 264:46:@33293.4]
  wire  _T_82; // @[Controllers.scala 264:62:@33294.4]
  wire  _T_100; // @[package.scala 100:49:@33312.4]
  reg  _T_103; // @[package.scala 48:56:@33313.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@33336.4]
  wire  _T_124; // @[package.scala 96:25:@33348.4 package.scala 96:25:@33349.4]
  wire  _T_126; // @[package.scala 100:49:@33350.4]
  reg  _T_129; // @[package.scala 48:56:@33351.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@33373.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@33375.4]
  reg  _T_153; // @[package.scala 48:56:@33376.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@33378.4]
  wire  _T_156; // @[Controllers.scala 292:61:@33379.4]
  wire  _T_157; // @[Controllers.scala 292:24:@33380.4]
  SRFF active ( // @[Controllers.scala 261:22:@33284.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@33287.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33321.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33343.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@33355.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@33363.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@33292.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@33293.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@33294.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@33312.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@33336.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33348.4 package.scala 96:25:@33349.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@33350.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@33375.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@33378.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@33379.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@33380.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@33354.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@33382.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@33339.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@33342.4]
  assign active_clock = clock; // @[:@33285.4]
  assign active_reset = reset; // @[:@33286.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@33297.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@33301.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@33302.4]
  assign done_clock = clock; // @[:@33288.4]
  assign done_reset = reset; // @[:@33289.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@33317.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@33310.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@33311.4]
  assign RetimeWrapper_clock = clock; // @[:@33322.4]
  assign RetimeWrapper_reset = reset; // @[:@33323.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33325.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@33324.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33344.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33345.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33347.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@33346.4]
  assign RetimeWrapper_2_clock = clock; // @[:@33356.4]
  assign RetimeWrapper_2_reset = reset; // @[:@33357.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@33359.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@33358.4]
  assign RetimeWrapper_3_clock = clock; // @[:@33364.4]
  assign RetimeWrapper_3_reset = reset; // @[:@33365.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@33367.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@33366.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1( // @[:@33457.2]
  output  io_in_x344_ready, // @[:@33460.4]
  input   io_sigsIn_datapathEn // @[:@33460.4]
);
  assign io_in_x344_ready = io_sigsIn_datapathEn; // @[sm_x362_inr_UnitPipe.scala 57:18:@33472.4]
endmodule
module x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1( // @[:@33475.2]
  input         clock, // @[:@33476.4]
  input         reset, // @[:@33477.4]
  output        io_in_x344_ready, // @[:@33478.4]
  input         io_in_x344_valid, // @[:@33478.4]
  output [20:0] io_in_x196_outbuf_0_rPort_0_ofs_0, // @[:@33478.4]
  output        io_in_x196_outbuf_0_rPort_0_en_0, // @[:@33478.4]
  output        io_in_x196_outbuf_0_rPort_0_backpressure, // @[:@33478.4]
  input  [31:0] io_in_x196_outbuf_0_rPort_0_output_0, // @[:@33478.4]
  input  [63:0] io_in_x192_outdram_number, // @[:@33478.4]
  input         io_in_x343_ready, // @[:@33478.4]
  output        io_in_x343_valid, // @[:@33478.4]
  output [31:0] io_in_x343_bits_wdata_0, // @[:@33478.4]
  output        io_in_x343_bits_wstrb, // @[:@33478.4]
  input         io_in_x342_ready, // @[:@33478.4]
  output        io_in_x342_valid, // @[:@33478.4]
  output [63:0] io_in_x342_bits_addr, // @[:@33478.4]
  output [31:0] io_in_x342_bits_size, // @[:@33478.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@33478.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@33478.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@33478.4]
  input         io_sigsIn_smChildAcks_0, // @[:@33478.4]
  input         io_sigsIn_smChildAcks_1, // @[:@33478.4]
  input         io_sigsIn_smChildAcks_2, // @[:@33478.4]
  output        io_sigsOut_smDoneIn_0, // @[:@33478.4]
  output        io_sigsOut_smDoneIn_1, // @[:@33478.4]
  output        io_sigsOut_smDoneIn_2, // @[:@33478.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@33478.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@33478.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@33478.4]
  input         io_rr // @[:@33478.4]
);
  wire  x349_inr_UnitPipe_sm_clock; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_reset; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_enable; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_done; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_doneLatch; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_ctrDone; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_datapathEn; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_ctrInc; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_parentAck; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  x349_inr_UnitPipe_sm_io_backpressure; // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33602.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33610.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33610.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33610.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33610.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33610.4]
  wire [63:0] x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x192_outdram_number; // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
  wire  x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_valid; // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
  wire [63:0] x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_bits_addr; // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
  wire [31:0] x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_bits_size; // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
  wire  x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
  wire  x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
  wire  x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_rr; // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
  wire  x351_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@33708.4]
  wire  x351_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@33708.4]
  wire  x351_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@33708.4]
  wire  x351_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@33708.4]
  wire [22:0] x351_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@33708.4]
  wire  x351_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@33708.4]
  wire  x351_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@33708.4]
  wire  x358_inr_Foreach_sm_clock; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_reset; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_enable; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_done; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_doneLatch; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_ctrDone; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_datapathEn; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_ctrInc; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_ctrRst; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_parentAck; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_backpressure; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  x358_inr_Foreach_sm_io_break; // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@33789.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@33789.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@33789.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@33789.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@33789.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@33829.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@33829.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@33829.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@33829.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@33829.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@33837.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@33837.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@33837.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@33837.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@33837.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_clock; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_reset; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire [20:0] x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_en_0; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire [31:0] x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_output_0; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_valid; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire [31:0] x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_bits_wdata_0; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_bits_wstrb; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire [31:0] x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_rr; // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
  wire  x362_inr_UnitPipe_sm_clock; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_reset; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_io_enable; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_io_done; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_io_doneLatch; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_io_ctrDone; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_io_datapathEn; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_io_ctrInc; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  x362_inr_UnitPipe_sm_io_parentAck; // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@34049.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@34049.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@34049.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@34049.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@34049.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@34057.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@34057.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@34057.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@34057.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@34057.4]
  wire  x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1_io_in_x344_ready; // @[sm_x362_inr_UnitPipe.scala 60:24:@34087.4]
  wire  x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x362_inr_UnitPipe.scala 60:24:@34087.4]
  wire  _T_359; // @[package.scala 100:49:@33573.4]
  reg  _T_362; // @[package.scala 48:56:@33574.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@33607.4 package.scala 96:25:@33608.4]
  wire  _T_381; // @[package.scala 96:25:@33615.4 package.scala 96:25:@33616.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@33618.4]
  wire  _T_454; // @[package.scala 96:25:@33794.4 package.scala 96:25:@33795.4]
  wire  _T_468; // @[package.scala 96:25:@33834.4 package.scala 96:25:@33835.4]
  wire  _T_474; // @[package.scala 96:25:@33842.4 package.scala 96:25:@33843.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@33845.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@33854.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@33855.4]
  wire  _T_547; // @[package.scala 100:49:@34020.4]
  reg  _T_550; // @[package.scala 48:56:@34021.4]
  reg [31:0] _RAND_1;
  wire  x362_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x363_outr_UnitPipe.scala 101:55:@34027.4]
  wire  _T_563; // @[package.scala 96:25:@34054.4 package.scala 96:25:@34055.4]
  wire  _T_569; // @[package.scala 96:25:@34062.4 package.scala 96:25:@34063.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@34065.4]
  wire  x362_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@34066.4]
  x349_inr_UnitPipe_sm x349_inr_UnitPipe_sm ( // @[sm_x349_inr_UnitPipe.scala 33:18:@33545.4]
    .clock(x349_inr_UnitPipe_sm_clock),
    .reset(x349_inr_UnitPipe_sm_reset),
    .io_enable(x349_inr_UnitPipe_sm_io_enable),
    .io_done(x349_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x349_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x349_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x349_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x349_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x349_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x349_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33602.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33610.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1 x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1 ( // @[sm_x349_inr_UnitPipe.scala 69:24:@33640.4]
    .io_in_x192_outdram_number(x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x192_outdram_number),
    .io_in_x342_valid(x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_valid),
    .io_in_x342_bits_addr(x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_bits_addr),
    .io_in_x342_bits_size(x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_bits_size),
    .io_sigsIn_backpressure(x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_rr)
  );
  x351_ctrchain x351_ctrchain ( // @[SpatialBlocks.scala 37:22:@33708.4]
    .clock(x351_ctrchain_clock),
    .reset(x351_ctrchain_reset),
    .io_input_reset(x351_ctrchain_io_input_reset),
    .io_input_enable(x351_ctrchain_io_input_enable),
    .io_output_counts_0(x351_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x351_ctrchain_io_output_oobs_0),
    .io_output_done(x351_ctrchain_io_output_done)
  );
  x358_inr_Foreach_sm x358_inr_Foreach_sm ( // @[sm_x358_inr_Foreach.scala 33:18:@33761.4]
    .clock(x358_inr_Foreach_sm_clock),
    .reset(x358_inr_Foreach_sm_reset),
    .io_enable(x358_inr_Foreach_sm_io_enable),
    .io_done(x358_inr_Foreach_sm_io_done),
    .io_doneLatch(x358_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x358_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x358_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x358_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x358_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x358_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x358_inr_Foreach_sm_io_backpressure),
    .io_break(x358_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@33789.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@33829.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@33837.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x358_inr_Foreach_kernelx358_inr_Foreach_concrete1 x358_inr_Foreach_kernelx358_inr_Foreach_concrete1 ( // @[sm_x358_inr_Foreach.scala 78:24:@33872.4]
    .clock(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_clock),
    .reset(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_reset),
    .io_in_x196_outbuf_0_rPort_0_ofs_0(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0),
    .io_in_x196_outbuf_0_rPort_0_en_0(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_en_0),
    .io_in_x196_outbuf_0_rPort_0_backpressure(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure),
    .io_in_x196_outbuf_0_rPort_0_output_0(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_output_0),
    .io_in_x343_valid(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_valid),
    .io_in_x343_bits_wdata_0(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_bits_wdata_0),
    .io_in_x343_bits_wstrb(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_bits_wstrb),
    .io_sigsIn_backpressure(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_rr)
  );
  x362_inr_UnitPipe_sm x362_inr_UnitPipe_sm ( // @[sm_x362_inr_UnitPipe.scala 32:18:@33992.4]
    .clock(x362_inr_UnitPipe_sm_clock),
    .reset(x362_inr_UnitPipe_sm_reset),
    .io_enable(x362_inr_UnitPipe_sm_io_enable),
    .io_done(x362_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x362_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x362_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x362_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x362_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x362_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@34049.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@34057.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1 x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1 ( // @[sm_x362_inr_UnitPipe.scala 60:24:@34087.4]
    .io_in_x344_ready(x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1_io_in_x344_ready),
    .io_sigsIn_datapathEn(x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x349_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33573.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@33607.4 package.scala 96:25:@33608.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33615.4 package.scala 96:25:@33616.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@33618.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@33794.4 package.scala 96:25:@33795.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@33834.4 package.scala 96:25:@33835.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@33842.4 package.scala 96:25:@33843.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@33845.4]
  assign _T_479 = x358_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@33854.4]
  assign _T_480 = ~ x358_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@33855.4]
  assign _T_547 = x362_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@34020.4]
  assign x362_inr_UnitPipe_sigsIn_forwardpressure = io_in_x344_valid | x362_inr_UnitPipe_sm_io_doneLatch; // @[sm_x363_outr_UnitPipe.scala 101:55:@34027.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@34054.4 package.scala 96:25:@34055.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@34062.4 package.scala 96:25:@34063.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@34065.4]
  assign x362_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@34066.4]
  assign io_in_x344_ready = x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1_io_in_x344_ready; // @[sm_x362_inr_UnitPipe.scala 46:23:@34123.4]
  assign io_in_x196_outbuf_0_rPort_0_ofs_0 = x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@33923.4]
  assign io_in_x196_outbuf_0_rPort_0_en_0 = x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@33922.4]
  assign io_in_x196_outbuf_0_rPort_0_backpressure = x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@33921.4]
  assign io_in_x343_valid = x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_valid; // @[sm_x358_inr_Foreach.scala 50:23:@33927.4]
  assign io_in_x343_bits_wdata_0 = x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_bits_wdata_0; // @[sm_x358_inr_Foreach.scala 50:23:@33926.4]
  assign io_in_x343_bits_wstrb = x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x343_bits_wstrb; // @[sm_x358_inr_Foreach.scala 50:23:@33925.4]
  assign io_in_x342_valid = x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_valid; // @[sm_x349_inr_UnitPipe.scala 50:23:@33679.4]
  assign io_in_x342_bits_addr = x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_bits_addr; // @[sm_x349_inr_UnitPipe.scala 50:23:@33678.4]
  assign io_in_x342_bits_size = x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x342_bits_size; // @[sm_x349_inr_UnitPipe.scala 50:23:@33677.4]
  assign io_sigsOut_smDoneIn_0 = x349_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33625.4]
  assign io_sigsOut_smDoneIn_1 = x358_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@33852.4]
  assign io_sigsOut_smDoneIn_2 = x362_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@34072.4]
  assign io_sigsOut_smCtrCopyDone_0 = x349_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@33639.4]
  assign io_sigsOut_smCtrCopyDone_1 = x358_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@33871.4]
  assign io_sigsOut_smCtrCopyDone_2 = x362_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@34086.4]
  assign x349_inr_UnitPipe_sm_clock = clock; // @[:@33546.4]
  assign x349_inr_UnitPipe_sm_reset = reset; // @[:@33547.4]
  assign x349_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@33622.4]
  assign x349_inr_UnitPipe_sm_io_ctrDone = x349_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x363_outr_UnitPipe.scala 77:39:@33577.4]
  assign x349_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@33624.4]
  assign x349_inr_UnitPipe_sm_io_backpressure = io_in_x342_ready | x349_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@33596.4]
  assign RetimeWrapper_clock = clock; // @[:@33603.4]
  assign RetimeWrapper_reset = reset; // @[:@33604.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33606.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@33605.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33611.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33612.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33614.4]
  assign RetimeWrapper_1_io_in = x349_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33613.4]
  assign x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_in_x192_outdram_number = io_in_x192_outdram_number; // @[sm_x349_inr_UnitPipe.scala 49:31:@33676.4]
  assign x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x342_ready | x349_inr_UnitPipe_sm_io_doneLatch; // @[sm_x349_inr_UnitPipe.scala 74:22:@33695.4]
  assign x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x349_inr_UnitPipe_sm_io_datapathEn; // @[sm_x349_inr_UnitPipe.scala 74:22:@33693.4]
  assign x349_inr_UnitPipe_kernelx349_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x349_inr_UnitPipe.scala 73:18:@33681.4]
  assign x351_ctrchain_clock = clock; // @[:@33709.4]
  assign x351_ctrchain_reset = reset; // @[:@33710.4]
  assign x351_ctrchain_io_input_reset = x358_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@33870.4]
  assign x351_ctrchain_io_input_enable = x358_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@33822.4 SpatialBlocks.scala 159:42:@33869.4]
  assign x358_inr_Foreach_sm_clock = clock; // @[:@33762.4]
  assign x358_inr_Foreach_sm_reset = reset; // @[:@33763.4]
  assign x358_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@33849.4]
  assign x358_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x363_outr_UnitPipe.scala 90:38:@33797.4]
  assign x358_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@33851.4]
  assign x358_inr_Foreach_sm_io_backpressure = io_in_x343_ready | x358_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@33823.4]
  assign x358_inr_Foreach_sm_io_break = 1'h0; // @[sm_x363_outr_UnitPipe.scala 94:36:@33803.4]
  assign RetimeWrapper_2_clock = clock; // @[:@33790.4]
  assign RetimeWrapper_2_reset = reset; // @[:@33791.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@33793.4]
  assign RetimeWrapper_2_io_in = x351_ctrchain_io_output_done; // @[package.scala 94:16:@33792.4]
  assign RetimeWrapper_3_clock = clock; // @[:@33830.4]
  assign RetimeWrapper_3_reset = reset; // @[:@33831.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@33833.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@33832.4]
  assign RetimeWrapper_4_clock = clock; // @[:@33838.4]
  assign RetimeWrapper_4_reset = reset; // @[:@33839.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@33841.4]
  assign RetimeWrapper_4_io_in = x358_inr_Foreach_sm_io_done; // @[package.scala 94:16:@33840.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_clock = clock; // @[:@33873.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_reset = reset; // @[:@33874.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_in_x196_outbuf_0_rPort_0_output_0 = io_in_x196_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@33920.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x343_ready | x358_inr_Foreach_sm_io_doneLatch; // @[sm_x358_inr_Foreach.scala 83:22:@33943.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x358_inr_Foreach.scala 83:22:@33941.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_break = x358_inr_Foreach_sm_io_break; // @[sm_x358_inr_Foreach.scala 83:22:@33939.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x351_ctrchain_io_output_counts_0[22]}},x351_ctrchain_io_output_counts_0}; // @[sm_x358_inr_Foreach.scala 83:22:@33934.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x351_ctrchain_io_output_oobs_0; // @[sm_x358_inr_Foreach.scala 83:22:@33933.4]
  assign x358_inr_Foreach_kernelx358_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x358_inr_Foreach.scala 82:18:@33929.4]
  assign x362_inr_UnitPipe_sm_clock = clock; // @[:@33993.4]
  assign x362_inr_UnitPipe_sm_reset = reset; // @[:@33994.4]
  assign x362_inr_UnitPipe_sm_io_enable = x362_inr_UnitPipe_sigsIn_baseEn & x362_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@34069.4]
  assign x362_inr_UnitPipe_sm_io_ctrDone = x362_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x363_outr_UnitPipe.scala 99:39:@34024.4]
  assign x362_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@34071.4]
  assign RetimeWrapper_5_clock = clock; // @[:@34050.4]
  assign RetimeWrapper_5_reset = reset; // @[:@34051.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@34053.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@34052.4]
  assign RetimeWrapper_6_clock = clock; // @[:@34058.4]
  assign RetimeWrapper_6_reset = reset; // @[:@34059.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@34061.4]
  assign RetimeWrapper_6_io_in = x362_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@34060.4]
  assign x362_inr_UnitPipe_kernelx362_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x362_inr_UnitPipe_sm_io_datapathEn; // @[sm_x362_inr_UnitPipe.scala 65:22:@34136.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x475_kernelx475_concrete1( // @[:@34152.2]
  input          clock, // @[:@34153.4]
  input          reset, // @[:@34154.4]
  output         io_in_x344_ready, // @[:@34155.4]
  input          io_in_x344_valid, // @[:@34155.4]
  output [20:0]  io_in_x196_outbuf_0_rPort_0_ofs_0, // @[:@34155.4]
  output         io_in_x196_outbuf_0_rPort_0_en_0, // @[:@34155.4]
  output         io_in_x196_outbuf_0_rPort_0_backpressure, // @[:@34155.4]
  input  [31:0]  io_in_x196_outbuf_0_rPort_0_output_0, // @[:@34155.4]
  input  [63:0]  io_in_x192_outdram_number, // @[:@34155.4]
  input          io_in_x343_ready, // @[:@34155.4]
  output         io_in_x343_valid, // @[:@34155.4]
  output [31:0]  io_in_x343_bits_wdata_0, // @[:@34155.4]
  output         io_in_x343_bits_wstrb, // @[:@34155.4]
  input          io_in_x342_ready, // @[:@34155.4]
  output         io_in_x342_valid, // @[:@34155.4]
  output [63:0]  io_in_x342_bits_addr, // @[:@34155.4]
  output [31:0]  io_in_x342_bits_size, // @[:@34155.4]
  input          io_in_x194_TVALID, // @[:@34155.4]
  output         io_in_x194_TREADY, // @[:@34155.4]
  input  [255:0] io_in_x194_TDATA, // @[:@34155.4]
  input  [7:0]   io_in_x194_TID, // @[:@34155.4]
  input  [7:0]   io_in_x194_TDEST, // @[:@34155.4]
  output         io_in_x195_TVALID, // @[:@34155.4]
  input          io_in_x195_TREADY, // @[:@34155.4]
  output [255:0] io_in_x195_TDATA, // @[:@34155.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@34155.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@34155.4]
  input          io_sigsIn_smChildAcks_0, // @[:@34155.4]
  input          io_sigsIn_smChildAcks_1, // @[:@34155.4]
  output         io_sigsOut_smDoneIn_0, // @[:@34155.4]
  output         io_sigsOut_smDoneIn_1, // @[:@34155.4]
  input          io_rr // @[:@34155.4]
);
  wire  x341_outr_UnitPipe_sm_clock; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_reset; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_enable; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_done; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_parentAck; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_childAck_0; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_childAck_1; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  x341_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34290.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34290.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34290.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34290.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34290.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34298.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34298.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34298.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34298.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34298.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_clock; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_reset; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TVALID; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TREADY; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire [255:0] x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TDATA; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire [7:0] x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TID; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire [7:0] x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TDEST; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TVALID; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TREADY; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire [255:0] x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TDATA; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_rr; // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
  wire  x363_outr_UnitPipe_sm_clock; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_reset; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_enable; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_done; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_parentAck; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_childAck_0; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_childAck_1; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_childAck_2; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  x363_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@34579.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@34579.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@34579.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@34579.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@34579.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@34587.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@34587.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@34587.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@34587.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@34587.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_clock; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_reset; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x344_ready; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x344_valid; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire [20:0] x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_en_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire [31:0] x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_output_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire [63:0] x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x192_outdram_number; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_ready; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_valid; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire [31:0] x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_bits_wdata_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_bits_wstrb; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_ready; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_valid; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire [63:0] x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_bits_addr; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire [31:0] x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_bits_size; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_rr; // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
  wire  _T_408; // @[package.scala 96:25:@34295.4 package.scala 96:25:@34296.4]
  wire  _T_414; // @[package.scala 96:25:@34303.4 package.scala 96:25:@34304.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@34306.4]
  wire  _T_508; // @[package.scala 96:25:@34584.4 package.scala 96:25:@34585.4]
  wire  _T_514; // @[package.scala 96:25:@34592.4 package.scala 96:25:@34593.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@34595.4]
  x341_outr_UnitPipe_sm x341_outr_UnitPipe_sm ( // @[sm_x341_outr_UnitPipe.scala 32:18:@34228.4]
    .clock(x341_outr_UnitPipe_sm_clock),
    .reset(x341_outr_UnitPipe_sm_reset),
    .io_enable(x341_outr_UnitPipe_sm_io_enable),
    .io_done(x341_outr_UnitPipe_sm_io_done),
    .io_parentAck(x341_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x341_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x341_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x341_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x341_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x341_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x341_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x341_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x341_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34290.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34298.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1 x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1 ( // @[sm_x341_outr_UnitPipe.scala 87:24:@34329.4]
    .clock(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_clock),
    .reset(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_reset),
    .io_in_x194_TVALID(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TVALID),
    .io_in_x194_TREADY(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TREADY),
    .io_in_x194_TDATA(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TDATA),
    .io_in_x194_TID(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TID),
    .io_in_x194_TDEST(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TDEST),
    .io_in_x195_TVALID(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TVALID),
    .io_in_x195_TREADY(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TREADY),
    .io_in_x195_TDATA(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TDATA),
    .io_sigsIn_smEnableOuts_0(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_rr)
  );
  x363_outr_UnitPipe_sm x363_outr_UnitPipe_sm ( // @[sm_x363_outr_UnitPipe.scala 36:18:@34507.4]
    .clock(x363_outr_UnitPipe_sm_clock),
    .reset(x363_outr_UnitPipe_sm_reset),
    .io_enable(x363_outr_UnitPipe_sm_io_enable),
    .io_done(x363_outr_UnitPipe_sm_io_done),
    .io_parentAck(x363_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x363_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x363_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x363_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x363_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x363_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x363_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x363_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x363_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x363_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x363_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x363_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x363_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@34579.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@34587.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1 x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1 ( // @[sm_x363_outr_UnitPipe.scala 108:24:@34619.4]
    .clock(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_clock),
    .reset(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_reset),
    .io_in_x344_ready(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x344_ready),
    .io_in_x344_valid(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x344_valid),
    .io_in_x196_outbuf_0_rPort_0_ofs_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0),
    .io_in_x196_outbuf_0_rPort_0_en_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_en_0),
    .io_in_x196_outbuf_0_rPort_0_backpressure(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure),
    .io_in_x196_outbuf_0_rPort_0_output_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_output_0),
    .io_in_x192_outdram_number(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x192_outdram_number),
    .io_in_x343_ready(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_ready),
    .io_in_x343_valid(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_valid),
    .io_in_x343_bits_wdata_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_bits_wdata_0),
    .io_in_x343_bits_wstrb(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_bits_wstrb),
    .io_in_x342_ready(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_ready),
    .io_in_x342_valid(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_valid),
    .io_in_x342_bits_addr(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_bits_addr),
    .io_in_x342_bits_size(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_bits_size),
    .io_sigsIn_smEnableOuts_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@34295.4 package.scala 96:25:@34296.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@34303.4 package.scala 96:25:@34304.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@34306.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@34584.4 package.scala 96:25:@34585.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@34592.4 package.scala 96:25:@34593.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@34595.4]
  assign io_in_x344_ready = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x344_ready; // @[sm_x363_outr_UnitPipe.scala 58:23:@34701.4]
  assign io_in_x196_outbuf_0_rPort_0_ofs_0 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@34705.4]
  assign io_in_x196_outbuf_0_rPort_0_en_0 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@34704.4]
  assign io_in_x196_outbuf_0_rPort_0_backpressure = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@34703.4]
  assign io_in_x343_valid = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_valid; // @[sm_x363_outr_UnitPipe.scala 61:23:@34710.4]
  assign io_in_x343_bits_wdata_0 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_bits_wdata_0; // @[sm_x363_outr_UnitPipe.scala 61:23:@34709.4]
  assign io_in_x343_bits_wstrb = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_bits_wstrb; // @[sm_x363_outr_UnitPipe.scala 61:23:@34708.4]
  assign io_in_x342_valid = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_valid; // @[sm_x363_outr_UnitPipe.scala 62:23:@34714.4]
  assign io_in_x342_bits_addr = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_bits_addr; // @[sm_x363_outr_UnitPipe.scala 62:23:@34713.4]
  assign io_in_x342_bits_size = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_bits_size; // @[sm_x363_outr_UnitPipe.scala 62:23:@34712.4]
  assign io_in_x194_TREADY = x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TREADY; // @[sm_x341_outr_UnitPipe.scala 48:23:@34397.4]
  assign io_in_x195_TVALID = x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TVALID; // @[sm_x341_outr_UnitPipe.scala 49:23:@34407.4]
  assign io_in_x195_TDATA = x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TDATA; // @[sm_x341_outr_UnitPipe.scala 49:23:@34405.4]
  assign io_sigsOut_smDoneIn_0 = x341_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@34313.4]
  assign io_sigsOut_smDoneIn_1 = x363_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@34602.4]
  assign x341_outr_UnitPipe_sm_clock = clock; // @[:@34229.4]
  assign x341_outr_UnitPipe_sm_reset = reset; // @[:@34230.4]
  assign x341_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@34310.4]
  assign x341_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@34312.4]
  assign x341_outr_UnitPipe_sm_io_doneIn_0 = x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@34280.4]
  assign x341_outr_UnitPipe_sm_io_doneIn_1 = x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@34281.4]
  assign x341_outr_UnitPipe_sm_io_ctrCopyDone_0 = x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@34327.4]
  assign x341_outr_UnitPipe_sm_io_ctrCopyDone_1 = x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@34328.4]
  assign RetimeWrapper_clock = clock; // @[:@34291.4]
  assign RetimeWrapper_reset = reset; // @[:@34292.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34294.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@34293.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34299.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34300.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34302.4]
  assign RetimeWrapper_1_io_in = x341_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@34301.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_clock = clock; // @[:@34330.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_reset = reset; // @[:@34331.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TVALID = io_in_x194_TVALID; // @[sm_x341_outr_UnitPipe.scala 48:23:@34398.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TDATA = io_in_x194_TDATA; // @[sm_x341_outr_UnitPipe.scala 48:23:@34396.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TID = io_in_x194_TID; // @[sm_x341_outr_UnitPipe.scala 48:23:@34392.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x194_TDEST = io_in_x194_TDEST; // @[sm_x341_outr_UnitPipe.scala 48:23:@34391.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_in_x195_TREADY = io_in_x195_TREADY; // @[sm_x341_outr_UnitPipe.scala 49:23:@34406.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x341_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x341_outr_UnitPipe.scala 92:22:@34423.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x341_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x341_outr_UnitPipe.scala 92:22:@34424.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x341_outr_UnitPipe_sm_io_childAck_0; // @[sm_x341_outr_UnitPipe.scala 92:22:@34419.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x341_outr_UnitPipe_sm_io_childAck_1; // @[sm_x341_outr_UnitPipe.scala 92:22:@34420.4]
  assign x341_outr_UnitPipe_kernelx341_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x341_outr_UnitPipe.scala 91:18:@34408.4]
  assign x363_outr_UnitPipe_sm_clock = clock; // @[:@34508.4]
  assign x363_outr_UnitPipe_sm_reset = reset; // @[:@34509.4]
  assign x363_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@34599.4]
  assign x363_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@34601.4]
  assign x363_outr_UnitPipe_sm_io_doneIn_0 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@34567.4]
  assign x363_outr_UnitPipe_sm_io_doneIn_1 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@34568.4]
  assign x363_outr_UnitPipe_sm_io_doneIn_2 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@34569.4]
  assign x363_outr_UnitPipe_sm_io_ctrCopyDone_0 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@34616.4]
  assign x363_outr_UnitPipe_sm_io_ctrCopyDone_1 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@34617.4]
  assign x363_outr_UnitPipe_sm_io_ctrCopyDone_2 = x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@34618.4]
  assign RetimeWrapper_2_clock = clock; // @[:@34580.4]
  assign RetimeWrapper_2_reset = reset; // @[:@34581.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@34583.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@34582.4]
  assign RetimeWrapper_3_clock = clock; // @[:@34588.4]
  assign RetimeWrapper_3_reset = reset; // @[:@34589.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@34591.4]
  assign RetimeWrapper_3_io_in = x363_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@34590.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_clock = clock; // @[:@34620.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_reset = reset; // @[:@34621.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x344_valid = io_in_x344_valid; // @[sm_x363_outr_UnitPipe.scala 58:23:@34700.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x196_outbuf_0_rPort_0_output_0 = io_in_x196_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@34702.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x192_outdram_number = io_in_x192_outdram_number; // @[sm_x363_outr_UnitPipe.scala 60:31:@34707.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x343_ready = io_in_x343_ready; // @[sm_x363_outr_UnitPipe.scala 61:23:@34711.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_in_x342_ready = io_in_x342_ready; // @[sm_x363_outr_UnitPipe.scala 62:23:@34715.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x363_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x363_outr_UnitPipe.scala 113:22:@34738.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x363_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x363_outr_UnitPipe.scala 113:22:@34739.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x363_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x363_outr_UnitPipe.scala 113:22:@34740.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x363_outr_UnitPipe_sm_io_childAck_0; // @[sm_x363_outr_UnitPipe.scala 113:22:@34732.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x363_outr_UnitPipe_sm_io_childAck_1; // @[sm_x363_outr_UnitPipe.scala 113:22:@34733.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x363_outr_UnitPipe_sm_io_childAck_2; // @[sm_x363_outr_UnitPipe.scala 113:22:@34734.4]
  assign x363_outr_UnitPipe_kernelx363_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x363_outr_UnitPipe.scala 112:18:@34716.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@34768.2]
  input          clock, // @[:@34769.4]
  input          reset, // @[:@34770.4]
  output         io_in_x344_ready, // @[:@34771.4]
  input          io_in_x344_valid, // @[:@34771.4]
  input  [63:0]  io_in_x192_outdram_number, // @[:@34771.4]
  input          io_in_x343_ready, // @[:@34771.4]
  output         io_in_x343_valid, // @[:@34771.4]
  output [31:0]  io_in_x343_bits_wdata_0, // @[:@34771.4]
  output         io_in_x343_bits_wstrb, // @[:@34771.4]
  input          io_in_x342_ready, // @[:@34771.4]
  output         io_in_x342_valid, // @[:@34771.4]
  output [63:0]  io_in_x342_bits_addr, // @[:@34771.4]
  output [31:0]  io_in_x342_bits_size, // @[:@34771.4]
  input          io_in_x194_TVALID, // @[:@34771.4]
  output         io_in_x194_TREADY, // @[:@34771.4]
  input  [255:0] io_in_x194_TDATA, // @[:@34771.4]
  input  [7:0]   io_in_x194_TID, // @[:@34771.4]
  input  [7:0]   io_in_x194_TDEST, // @[:@34771.4]
  output         io_in_x195_TVALID, // @[:@34771.4]
  input          io_in_x195_TREADY, // @[:@34771.4]
  output [255:0] io_in_x195_TDATA, // @[:@34771.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@34771.4]
  input          io_sigsIn_smChildAcks_0, // @[:@34771.4]
  output         io_sigsOut_smDoneIn_0, // @[:@34771.4]
  input          io_rr // @[:@34771.4]
);
  wire  x196_outbuf_0_clock; // @[m_x196_outbuf_0.scala 27:17:@34781.4]
  wire  x196_outbuf_0_reset; // @[m_x196_outbuf_0.scala 27:17:@34781.4]
  wire [20:0] x196_outbuf_0_io_rPort_0_ofs_0; // @[m_x196_outbuf_0.scala 27:17:@34781.4]
  wire  x196_outbuf_0_io_rPort_0_en_0; // @[m_x196_outbuf_0.scala 27:17:@34781.4]
  wire  x196_outbuf_0_io_rPort_0_backpressure; // @[m_x196_outbuf_0.scala 27:17:@34781.4]
  wire [31:0] x196_outbuf_0_io_rPort_0_output_0; // @[m_x196_outbuf_0.scala 27:17:@34781.4]
  wire  x475_sm_clock; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_reset; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_enable; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_done; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_ctrDone; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_ctrInc; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_parentAck; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_doneIn_0; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_doneIn_1; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_enableOut_0; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_enableOut_1; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_childAck_0; // @[sm_x475.scala 37:18:@34839.4]
  wire  x475_sm_io_childAck_1; // @[sm_x475.scala 37:18:@34839.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34914.4]
  wire  x475_kernelx475_concrete1_clock; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_reset; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x344_ready; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x344_valid; // @[sm_x475.scala 102:24:@34943.4]
  wire [20:0] x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_en_0; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure; // @[sm_x475.scala 102:24:@34943.4]
  wire [31:0] x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_output_0; // @[sm_x475.scala 102:24:@34943.4]
  wire [63:0] x475_kernelx475_concrete1_io_in_x192_outdram_number; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x343_ready; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x343_valid; // @[sm_x475.scala 102:24:@34943.4]
  wire [31:0] x475_kernelx475_concrete1_io_in_x343_bits_wdata_0; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x343_bits_wstrb; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x342_ready; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x342_valid; // @[sm_x475.scala 102:24:@34943.4]
  wire [63:0] x475_kernelx475_concrete1_io_in_x342_bits_addr; // @[sm_x475.scala 102:24:@34943.4]
  wire [31:0] x475_kernelx475_concrete1_io_in_x342_bits_size; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x194_TVALID; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x194_TREADY; // @[sm_x475.scala 102:24:@34943.4]
  wire [255:0] x475_kernelx475_concrete1_io_in_x194_TDATA; // @[sm_x475.scala 102:24:@34943.4]
  wire [7:0] x475_kernelx475_concrete1_io_in_x194_TID; // @[sm_x475.scala 102:24:@34943.4]
  wire [7:0] x475_kernelx475_concrete1_io_in_x194_TDEST; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x195_TVALID; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_in_x195_TREADY; // @[sm_x475.scala 102:24:@34943.4]
  wire [255:0] x475_kernelx475_concrete1_io_in_x195_TDATA; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x475.scala 102:24:@34943.4]
  wire  x475_kernelx475_concrete1_io_rr; // @[sm_x475.scala 102:24:@34943.4]
  wire  _T_266; // @[package.scala 100:49:@34872.4]
  reg  _T_269; // @[package.scala 48:56:@34873.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@34911.4 package.scala 96:25:@34912.4]
  wire  _T_289; // @[package.scala 96:25:@34919.4 package.scala 96:25:@34920.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@34922.4]
  x196_outbuf_0 x196_outbuf_0 ( // @[m_x196_outbuf_0.scala 27:17:@34781.4]
    .clock(x196_outbuf_0_clock),
    .reset(x196_outbuf_0_reset),
    .io_rPort_0_ofs_0(x196_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x196_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x196_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x196_outbuf_0_io_rPort_0_output_0)
  );
  x475_sm x475_sm ( // @[sm_x475.scala 37:18:@34839.4]
    .clock(x475_sm_clock),
    .reset(x475_sm_reset),
    .io_enable(x475_sm_io_enable),
    .io_done(x475_sm_io_done),
    .io_ctrDone(x475_sm_io_ctrDone),
    .io_ctrInc(x475_sm_io_ctrInc),
    .io_parentAck(x475_sm_io_parentAck),
    .io_doneIn_0(x475_sm_io_doneIn_0),
    .io_doneIn_1(x475_sm_io_doneIn_1),
    .io_enableOut_0(x475_sm_io_enableOut_0),
    .io_enableOut_1(x475_sm_io_enableOut_1),
    .io_childAck_0(x475_sm_io_childAck_0),
    .io_childAck_1(x475_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34906.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34914.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x475_kernelx475_concrete1 x475_kernelx475_concrete1 ( // @[sm_x475.scala 102:24:@34943.4]
    .clock(x475_kernelx475_concrete1_clock),
    .reset(x475_kernelx475_concrete1_reset),
    .io_in_x344_ready(x475_kernelx475_concrete1_io_in_x344_ready),
    .io_in_x344_valid(x475_kernelx475_concrete1_io_in_x344_valid),
    .io_in_x196_outbuf_0_rPort_0_ofs_0(x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0),
    .io_in_x196_outbuf_0_rPort_0_en_0(x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_en_0),
    .io_in_x196_outbuf_0_rPort_0_backpressure(x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure),
    .io_in_x196_outbuf_0_rPort_0_output_0(x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_output_0),
    .io_in_x192_outdram_number(x475_kernelx475_concrete1_io_in_x192_outdram_number),
    .io_in_x343_ready(x475_kernelx475_concrete1_io_in_x343_ready),
    .io_in_x343_valid(x475_kernelx475_concrete1_io_in_x343_valid),
    .io_in_x343_bits_wdata_0(x475_kernelx475_concrete1_io_in_x343_bits_wdata_0),
    .io_in_x343_bits_wstrb(x475_kernelx475_concrete1_io_in_x343_bits_wstrb),
    .io_in_x342_ready(x475_kernelx475_concrete1_io_in_x342_ready),
    .io_in_x342_valid(x475_kernelx475_concrete1_io_in_x342_valid),
    .io_in_x342_bits_addr(x475_kernelx475_concrete1_io_in_x342_bits_addr),
    .io_in_x342_bits_size(x475_kernelx475_concrete1_io_in_x342_bits_size),
    .io_in_x194_TVALID(x475_kernelx475_concrete1_io_in_x194_TVALID),
    .io_in_x194_TREADY(x475_kernelx475_concrete1_io_in_x194_TREADY),
    .io_in_x194_TDATA(x475_kernelx475_concrete1_io_in_x194_TDATA),
    .io_in_x194_TID(x475_kernelx475_concrete1_io_in_x194_TID),
    .io_in_x194_TDEST(x475_kernelx475_concrete1_io_in_x194_TDEST),
    .io_in_x195_TVALID(x475_kernelx475_concrete1_io_in_x195_TVALID),
    .io_in_x195_TREADY(x475_kernelx475_concrete1_io_in_x195_TREADY),
    .io_in_x195_TDATA(x475_kernelx475_concrete1_io_in_x195_TDATA),
    .io_sigsIn_smEnableOuts_0(x475_kernelx475_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x475_kernelx475_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x475_kernelx475_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x475_kernelx475_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x475_kernelx475_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x475_kernelx475_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x475_kernelx475_concrete1_io_rr)
  );
  assign _T_266 = x475_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@34872.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@34911.4 package.scala 96:25:@34912.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@34919.4 package.scala 96:25:@34920.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@34922.4]
  assign io_in_x344_ready = x475_kernelx475_concrete1_io_in_x344_ready; // @[sm_x475.scala 63:23:@35024.4]
  assign io_in_x343_valid = x475_kernelx475_concrete1_io_in_x343_valid; // @[sm_x475.scala 66:23:@35033.4]
  assign io_in_x343_bits_wdata_0 = x475_kernelx475_concrete1_io_in_x343_bits_wdata_0; // @[sm_x475.scala 66:23:@35032.4]
  assign io_in_x343_bits_wstrb = x475_kernelx475_concrete1_io_in_x343_bits_wstrb; // @[sm_x475.scala 66:23:@35031.4]
  assign io_in_x342_valid = x475_kernelx475_concrete1_io_in_x342_valid; // @[sm_x475.scala 67:23:@35037.4]
  assign io_in_x342_bits_addr = x475_kernelx475_concrete1_io_in_x342_bits_addr; // @[sm_x475.scala 67:23:@35036.4]
  assign io_in_x342_bits_size = x475_kernelx475_concrete1_io_in_x342_bits_size; // @[sm_x475.scala 67:23:@35035.4]
  assign io_in_x194_TREADY = x475_kernelx475_concrete1_io_in_x194_TREADY; // @[sm_x475.scala 68:23:@35046.4]
  assign io_in_x195_TVALID = x475_kernelx475_concrete1_io_in_x195_TVALID; // @[sm_x475.scala 69:23:@35056.4]
  assign io_in_x195_TDATA = x475_kernelx475_concrete1_io_in_x195_TDATA; // @[sm_x475.scala 69:23:@35054.4]
  assign io_sigsOut_smDoneIn_0 = x475_sm_io_done; // @[SpatialBlocks.scala 156:53:@34929.4]
  assign x196_outbuf_0_clock = clock; // @[:@34782.4]
  assign x196_outbuf_0_reset = reset; // @[:@34783.4]
  assign x196_outbuf_0_io_rPort_0_ofs_0 = x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@35028.4]
  assign x196_outbuf_0_io_rPort_0_en_0 = x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@35027.4]
  assign x196_outbuf_0_io_rPort_0_backpressure = x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@35026.4]
  assign x475_sm_clock = clock; // @[:@34840.4]
  assign x475_sm_reset = reset; // @[:@34841.4]
  assign x475_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@34926.4]
  assign x475_sm_io_ctrDone = x475_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@34876.4]
  assign x475_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@34928.4]
  assign x475_sm_io_doneIn_0 = x475_kernelx475_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@34896.4]
  assign x475_sm_io_doneIn_1 = x475_kernelx475_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@34897.4]
  assign RetimeWrapper_clock = clock; // @[:@34907.4]
  assign RetimeWrapper_reset = reset; // @[:@34908.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34910.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@34909.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34915.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34916.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34918.4]
  assign RetimeWrapper_1_io_in = x475_sm_io_done; // @[package.scala 94:16:@34917.4]
  assign x475_kernelx475_concrete1_clock = clock; // @[:@34944.4]
  assign x475_kernelx475_concrete1_reset = reset; // @[:@34945.4]
  assign x475_kernelx475_concrete1_io_in_x344_valid = io_in_x344_valid; // @[sm_x475.scala 63:23:@35023.4]
  assign x475_kernelx475_concrete1_io_in_x196_outbuf_0_rPort_0_output_0 = x196_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@35025.4]
  assign x475_kernelx475_concrete1_io_in_x192_outdram_number = io_in_x192_outdram_number; // @[sm_x475.scala 65:31:@35030.4]
  assign x475_kernelx475_concrete1_io_in_x343_ready = io_in_x343_ready; // @[sm_x475.scala 66:23:@35034.4]
  assign x475_kernelx475_concrete1_io_in_x342_ready = io_in_x342_ready; // @[sm_x475.scala 67:23:@35038.4]
  assign x475_kernelx475_concrete1_io_in_x194_TVALID = io_in_x194_TVALID; // @[sm_x475.scala 68:23:@35047.4]
  assign x475_kernelx475_concrete1_io_in_x194_TDATA = io_in_x194_TDATA; // @[sm_x475.scala 68:23:@35045.4]
  assign x475_kernelx475_concrete1_io_in_x194_TID = io_in_x194_TID; // @[sm_x475.scala 68:23:@35041.4]
  assign x475_kernelx475_concrete1_io_in_x194_TDEST = io_in_x194_TDEST; // @[sm_x475.scala 68:23:@35040.4]
  assign x475_kernelx475_concrete1_io_in_x195_TREADY = io_in_x195_TREADY; // @[sm_x475.scala 69:23:@35055.4]
  assign x475_kernelx475_concrete1_io_sigsIn_smEnableOuts_0 = x475_sm_io_enableOut_0; // @[sm_x475.scala 107:22:@35067.4]
  assign x475_kernelx475_concrete1_io_sigsIn_smEnableOuts_1 = x475_sm_io_enableOut_1; // @[sm_x475.scala 107:22:@35068.4]
  assign x475_kernelx475_concrete1_io_sigsIn_smChildAcks_0 = x475_sm_io_childAck_0; // @[sm_x475.scala 107:22:@35063.4]
  assign x475_kernelx475_concrete1_io_sigsIn_smChildAcks_1 = x475_sm_io_childAck_1; // @[sm_x475.scala 107:22:@35064.4]
  assign x475_kernelx475_concrete1_io_rr = io_rr; // @[sm_x475.scala 106:18:@35057.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@35090.2]
  input          clock, // @[:@35091.4]
  input          reset, // @[:@35092.4]
  input          io_enable, // @[:@35093.4]
  output         io_done, // @[:@35093.4]
  input          io_reset, // @[:@35093.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@35093.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@35093.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@35093.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@35093.4]
  output         io_memStreams_loads_0_data_ready, // @[:@35093.4]
  input          io_memStreams_loads_0_data_valid, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@35093.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@35093.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@35093.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@35093.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@35093.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@35093.4]
  input          io_memStreams_stores_0_data_ready, // @[:@35093.4]
  output         io_memStreams_stores_0_data_valid, // @[:@35093.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@35093.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@35093.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@35093.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@35093.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@35093.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@35093.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@35093.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@35093.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@35093.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@35093.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@35093.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@35093.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@35093.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@35093.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@35093.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@35093.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@35093.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@35093.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@35093.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@35093.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@35093.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@35093.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@35093.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@35093.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@35093.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@35093.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@35093.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@35093.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@35093.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@35093.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@35093.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@35093.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@35093.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@35093.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@35093.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@35093.4]
  output         io_heap_0_req_valid, // @[:@35093.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@35093.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@35093.4]
  input          io_heap_0_resp_valid, // @[:@35093.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@35093.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@35093.4]
  input  [63:0]  io_argIns_0, // @[:@35093.4]
  input  [63:0]  io_argIns_1, // @[:@35093.4]
  input          io_argOuts_0_port_ready, // @[:@35093.4]
  output         io_argOuts_0_port_valid, // @[:@35093.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@35093.4]
  input  [63:0]  io_argOuts_0_echo // @[:@35093.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@35241.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@35241.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@35241.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@35241.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@35259.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@35259.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@35259.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@35259.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@35259.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@35268.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@35268.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@35268.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@35268.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@35268.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@35268.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@35307.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@35339.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@35339.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@35339.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@35339.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@35339.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x344_ready; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x344_valid; // @[sm_RootController.scala 91:24:@35401.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x192_outdram_number; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x343_ready; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x343_valid; // @[sm_RootController.scala 91:24:@35401.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x343_bits_wdata_0; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x343_bits_wstrb; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x342_ready; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x342_valid; // @[sm_RootController.scala 91:24:@35401.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x342_bits_addr; // @[sm_RootController.scala 91:24:@35401.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x342_bits_size; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x194_TVALID; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x194_TREADY; // @[sm_RootController.scala 91:24:@35401.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x194_TDATA; // @[sm_RootController.scala 91:24:@35401.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x194_TID; // @[sm_RootController.scala 91:24:@35401.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x194_TDEST; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x195_TVALID; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_in_x195_TREADY; // @[sm_RootController.scala 91:24:@35401.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x195_TDATA; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@35401.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@35401.4]
  wire  _T_599; // @[package.scala 96:25:@35264.4 package.scala 96:25:@35265.4]
  wire  _T_664; // @[Main.scala 46:50:@35335.4]
  wire  _T_665; // @[Main.scala 46:59:@35336.4]
  wire  _T_677; // @[package.scala 100:49:@35356.4]
  reg  _T_680; // @[package.scala 48:56:@35357.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@35241.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@35259.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@35268.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@35307.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@35339.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@35401.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x344_ready(RootController_kernelRootController_concrete1_io_in_x344_ready),
    .io_in_x344_valid(RootController_kernelRootController_concrete1_io_in_x344_valid),
    .io_in_x192_outdram_number(RootController_kernelRootController_concrete1_io_in_x192_outdram_number),
    .io_in_x343_ready(RootController_kernelRootController_concrete1_io_in_x343_ready),
    .io_in_x343_valid(RootController_kernelRootController_concrete1_io_in_x343_valid),
    .io_in_x343_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x343_bits_wdata_0),
    .io_in_x343_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x343_bits_wstrb),
    .io_in_x342_ready(RootController_kernelRootController_concrete1_io_in_x342_ready),
    .io_in_x342_valid(RootController_kernelRootController_concrete1_io_in_x342_valid),
    .io_in_x342_bits_addr(RootController_kernelRootController_concrete1_io_in_x342_bits_addr),
    .io_in_x342_bits_size(RootController_kernelRootController_concrete1_io_in_x342_bits_size),
    .io_in_x194_TVALID(RootController_kernelRootController_concrete1_io_in_x194_TVALID),
    .io_in_x194_TREADY(RootController_kernelRootController_concrete1_io_in_x194_TREADY),
    .io_in_x194_TDATA(RootController_kernelRootController_concrete1_io_in_x194_TDATA),
    .io_in_x194_TID(RootController_kernelRootController_concrete1_io_in_x194_TID),
    .io_in_x194_TDEST(RootController_kernelRootController_concrete1_io_in_x194_TDEST),
    .io_in_x195_TVALID(RootController_kernelRootController_concrete1_io_in_x195_TVALID),
    .io_in_x195_TREADY(RootController_kernelRootController_concrete1_io_in_x195_TREADY),
    .io_in_x195_TDATA(RootController_kernelRootController_concrete1_io_in_x195_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@35264.4 package.scala 96:25:@35265.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@35335.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@35336.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@35356.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@35355.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x342_valid; // @[sm_RootController.scala 63:23:@35472.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x342_bits_addr; // @[sm_RootController.scala 63:23:@35471.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x342_bits_size; // @[sm_RootController.scala 63:23:@35470.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x343_valid; // @[sm_RootController.scala 62:23:@35468.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x343_bits_wdata_0; // @[sm_RootController.scala 62:23:@35467.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x343_bits_wstrb; // @[sm_RootController.scala 62:23:@35466.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x344_ready; // @[sm_RootController.scala 60:23:@35464.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x194_TREADY; // @[sm_RootController.scala 64:23:@35481.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x195_TVALID; // @[sm_RootController.scala 65:23:@35491.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x195_TDATA; // @[sm_RootController.scala 65:23:@35489.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 65:23:@35488.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 65:23:@35487.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 65:23:@35486.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 65:23:@35485.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 65:23:@35484.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 65:23:@35483.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@35242.4]
  assign SingleCounter_reset = reset; // @[:@35243.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@35257.4]
  assign RetimeWrapper_clock = clock; // @[:@35260.4]
  assign RetimeWrapper_reset = reset; // @[:@35261.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@35263.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@35262.4]
  assign SRFF_clock = clock; // @[:@35269.4]
  assign SRFF_reset = reset; // @[:@35270.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@35519.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@35353.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@35354.4]
  assign RootController_sm_clock = clock; // @[:@35308.4]
  assign RootController_sm_reset = reset; // @[:@35309.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@35352.4 SpatialBlocks.scala 140:18:@35386.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@35380.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@35360.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@35348.4 SpatialBlocks.scala 142:21:@35388.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@35377.4]
  assign RetimeWrapper_1_clock = clock; // @[:@35340.4]
  assign RetimeWrapper_1_reset = reset; // @[:@35341.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@35343.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@35342.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@35402.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@35403.4]
  assign RootController_kernelRootController_concrete1_io_in_x344_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 60:23:@35463.4]
  assign RootController_kernelRootController_concrete1_io_in_x192_outdram_number = io_argIns_1; // @[sm_RootController.scala 61:31:@35465.4]
  assign RootController_kernelRootController_concrete1_io_in_x343_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 62:23:@35469.4]
  assign RootController_kernelRootController_concrete1_io_in_x342_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 63:23:@35473.4]
  assign RootController_kernelRootController_concrete1_io_in_x194_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 64:23:@35482.4]
  assign RootController_kernelRootController_concrete1_io_in_x194_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 64:23:@35480.4]
  assign RootController_kernelRootController_concrete1_io_in_x194_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 64:23:@35476.4]
  assign RootController_kernelRootController_concrete1_io_in_x194_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 64:23:@35475.4]
  assign RootController_kernelRootController_concrete1_io_in_x195_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 65:23:@35490.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@35500.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@35498.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@35492.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@35521.2]
  input        clock, // @[:@35522.4]
  input        reset, // @[:@35523.4]
  input        io_enable, // @[:@35524.4]
  output [5:0] io_out, // @[:@35524.4]
  output [5:0] io_next // @[:@35524.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@35526.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@35527.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@35528.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@35533.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@35527.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@35528.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@35533.6]
  assign io_out = count; // @[Counter.scala 25:10:@35536.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@35537.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_13( // @[:@35573.2]
  input         clock, // @[:@35574.4]
  input         reset, // @[:@35575.4]
  input  [5:0]  io_raddr, // @[:@35576.4]
  input         io_wen, // @[:@35576.4]
  input  [5:0]  io_waddr, // @[:@35576.4]
  input  [63:0] io_wdata_addr, // @[:@35576.4]
  input  [31:0] io_wdata_size, // @[:@35576.4]
  output [63:0] io_rdata_addr, // @[:@35576.4]
  output [31:0] io_rdata_size // @[:@35576.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@35578.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@35578.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@35578.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@35578.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@35578.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@35578.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@35578.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@35578.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@35578.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@35592.4]
  wire  _T_20; // @[SRAM.scala 182:49:@35597.4]
  wire  _T_21; // @[SRAM.scala 182:37:@35598.4]
  reg  _T_24; // @[SRAM.scala 182:29:@35599.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@35602.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@35604.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@35578.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@35592.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@35597.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@35598.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@35604.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@35613.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@35612.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@35593.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@35594.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@35590.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@35596.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@35595.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@35591.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@35589.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@35588.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@35615.2]
  input         clock, // @[:@35616.4]
  input         reset, // @[:@35617.4]
  output        io_in_ready, // @[:@35618.4]
  input         io_in_valid, // @[:@35618.4]
  input  [63:0] io_in_bits_addr, // @[:@35618.4]
  input  [31:0] io_in_bits_size, // @[:@35618.4]
  input         io_out_ready, // @[:@35618.4]
  output        io_out_valid, // @[:@35618.4]
  output [63:0] io_out_bits_addr, // @[:@35618.4]
  output [31:0] io_out_bits_size // @[:@35618.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@36014.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@36014.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@36014.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@36014.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@36014.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@36024.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@36024.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@36024.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@36024.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@36024.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@36039.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@36039.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@36039.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@36039.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@36039.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@36039.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@36039.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@36039.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@36039.4]
  wire  writeEn; // @[FIFO.scala 30:29:@36012.4]
  wire  readEn; // @[FIFO.scala 31:29:@36013.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@36034.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@36035.4]
  wire  _T_824; // @[FIFO.scala 45:27:@36036.4]
  wire  empty; // @[FIFO.scala 45:24:@36037.4]
  wire  full; // @[FIFO.scala 46:23:@36038.4]
  wire  _T_827; // @[FIFO.scala 83:17:@36051.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@36052.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@36014.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@36024.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_13 SRAM ( // @[FIFO.scala 73:19:@36039.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@36012.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@36013.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@36035.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@36036.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@36037.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@36038.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@36051.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@36052.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@36058.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@36056.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@36049.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@36048.4]
  assign enqCounter_clock = clock; // @[:@36015.4]
  assign enqCounter_reset = reset; // @[:@36016.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@36022.4]
  assign deqCounter_clock = clock; // @[:@36025.4]
  assign deqCounter_reset = reset; // @[:@36026.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@36032.4]
  assign SRAM_clock = clock; // @[:@36040.4]
  assign SRAM_reset = reset; // @[:@36041.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@36043.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@36044.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@36045.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@36047.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@36046.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@36060.2]
  input        clock, // @[:@36061.4]
  input        reset, // @[:@36062.4]
  input        io_enable, // @[:@36063.4]
  output [3:0] io_out // @[:@36063.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@36065.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@36066.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@36067.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@36072.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@36066.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@36067.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@36072.6]
  assign io_out = count; // @[Counter.scala 25:10:@36075.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@36096.2]
  input        clock, // @[:@36097.4]
  input        reset, // @[:@36098.4]
  input        io_reset, // @[:@36099.4]
  input        io_enable, // @[:@36099.4]
  input  [1:0] io_stride, // @[:@36099.4]
  output [1:0] io_out, // @[:@36099.4]
  output [1:0] io_next // @[:@36099.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@36101.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@36102.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@36103.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@36108.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@36104.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@36102.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@36103.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@36108.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@36104.4]
  assign io_out = count; // @[Counter.scala 25:10:@36111.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@36112.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_14( // @[:@36148.2]
  input         clock, // @[:@36149.4]
  input         reset, // @[:@36150.4]
  input  [1:0]  io_raddr, // @[:@36151.4]
  input         io_wen, // @[:@36151.4]
  input  [1:0]  io_waddr, // @[:@36151.4]
  input  [31:0] io_wdata, // @[:@36151.4]
  output [31:0] io_rdata, // @[:@36151.4]
  input         io_backpressure // @[:@36151.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@36153.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@36153.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@36153.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@36153.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@36153.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@36153.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@36153.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@36153.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@36153.4]
  wire  _T_19; // @[SRAM.scala 182:49:@36171.4]
  wire  _T_20; // @[SRAM.scala 182:37:@36172.4]
  reg  _T_23; // @[SRAM.scala 182:29:@36173.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@36175.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@36153.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@36171.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@36172.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@36180.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@36167.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@36168.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@36165.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@36170.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@36169.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@36166.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@36164.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@36163.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@36182.2]
  input         clock, // @[:@36183.4]
  input         reset, // @[:@36184.4]
  output        io_in_ready, // @[:@36185.4]
  input         io_in_valid, // @[:@36185.4]
  input  [31:0] io_in_bits, // @[:@36185.4]
  input         io_out_ready, // @[:@36185.4]
  output        io_out_valid, // @[:@36185.4]
  output [31:0] io_out_bits // @[:@36185.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@36211.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@36211.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@36211.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@36211.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@36211.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@36211.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@36211.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@36221.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@36221.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@36221.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@36221.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@36221.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@36221.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@36221.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@36236.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@36236.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@36236.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@36236.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@36236.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@36236.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@36236.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@36236.4]
  wire  writeEn; // @[FIFO.scala 30:29:@36209.4]
  wire  readEn; // @[FIFO.scala 31:29:@36210.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@36231.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@36232.4]
  wire  _T_104; // @[FIFO.scala 45:27:@36233.4]
  wire  empty; // @[FIFO.scala 45:24:@36234.4]
  wire  full; // @[FIFO.scala 46:23:@36235.4]
  wire  _T_107; // @[FIFO.scala 83:17:@36246.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@36247.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@36211.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@36221.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_14 SRAM ( // @[FIFO.scala 73:19:@36236.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@36209.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@36210.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@36232.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@36233.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@36234.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@36235.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@36246.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@36247.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@36253.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@36251.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@36244.4]
  assign enqCounter_clock = clock; // @[:@36212.4]
  assign enqCounter_reset = reset; // @[:@36213.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@36219.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@36220.4]
  assign deqCounter_clock = clock; // @[:@36222.4]
  assign deqCounter_reset = reset; // @[:@36223.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@36229.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@36230.4]
  assign SRAM_clock = clock; // @[:@36237.4]
  assign SRAM_reset = reset; // @[:@36238.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@36240.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@36241.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@36242.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@36243.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@36245.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@38640.2]
  input         clock, // @[:@38641.4]
  input         reset, // @[:@38642.4]
  output        io_in_ready, // @[:@38643.4]
  input         io_in_valid, // @[:@38643.4]
  input  [31:0] io_in_bits_0, // @[:@38643.4]
  input         io_out_ready, // @[:@38643.4]
  output        io_out_valid, // @[:@38643.4]
  output [31:0] io_out_bits_0, // @[:@38643.4]
  output [31:0] io_out_bits_1, // @[:@38643.4]
  output [31:0] io_out_bits_2, // @[:@38643.4]
  output [31:0] io_out_bits_3, // @[:@38643.4]
  output [31:0] io_out_bits_4, // @[:@38643.4]
  output [31:0] io_out_bits_5, // @[:@38643.4]
  output [31:0] io_out_bits_6, // @[:@38643.4]
  output [31:0] io_out_bits_7, // @[:@38643.4]
  output [31:0] io_out_bits_8, // @[:@38643.4]
  output [31:0] io_out_bits_9, // @[:@38643.4]
  output [31:0] io_out_bits_10, // @[:@38643.4]
  output [31:0] io_out_bits_11, // @[:@38643.4]
  output [31:0] io_out_bits_12, // @[:@38643.4]
  output [31:0] io_out_bits_13, // @[:@38643.4]
  output [31:0] io_out_bits_14, // @[:@38643.4]
  output [31:0] io_out_bits_15 // @[:@38643.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@38647.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@38647.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@38647.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@38647.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@38658.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@38658.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@38658.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@38658.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@38671.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@38671.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@38671.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@38671.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@38671.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@38671.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@38671.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@38671.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@38706.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@38706.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@38706.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@38706.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@38706.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@38706.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@38706.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@38706.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@38741.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@38741.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@38741.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@38741.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@38741.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@38741.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@38741.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@38741.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@38776.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@38776.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@38776.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@38776.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@38776.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@38776.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@38776.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@38776.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@38811.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@38811.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@38811.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@38811.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@38811.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@38811.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@38811.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@38811.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@38846.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@38846.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@38846.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@38846.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@38846.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@38846.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@38846.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@38846.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@38881.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@38881.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@38881.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@38881.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@38881.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@38881.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@38881.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@38881.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@38916.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@38916.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@38916.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@38916.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@38916.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@38916.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@38916.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@38916.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@38951.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@38951.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@38951.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@38951.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@38951.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@38951.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@38951.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@38951.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@38986.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@38986.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@38986.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@38986.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@38986.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@38986.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@38986.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@38986.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@39021.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@39021.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@39021.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@39021.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@39021.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@39021.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@39021.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@39021.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@39056.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@39056.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@39056.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@39056.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@39056.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@39056.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@39056.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@39056.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@39091.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@39091.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@39091.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@39091.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@39091.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@39091.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@39091.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@39091.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@39126.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@39126.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@39126.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@39126.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@39126.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@39126.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@39126.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@39126.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@39161.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@39161.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@39161.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@39161.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@39161.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@39161.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@39161.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@39161.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@39196.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@39196.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@39196.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@39196.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@39196.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@39196.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@39196.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@39196.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@38646.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@38669.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@38696.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@38731.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@38766.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@38801.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@38836.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@38871.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@38906.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@38941.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@38976.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@39011.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@39046.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@39081.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@39116.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@39151.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@39186.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@39221.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39232.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39233.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39234.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39235.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39236.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39237.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39238.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39239.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39240.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39241.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39242.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39243.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39244.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39245.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39246.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@39263.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39247.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@39282.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@39283.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@39284.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@39285.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@39286.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@39287.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@39288.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@39289.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@39290.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@39291.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@39292.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@39293.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@39294.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@39295.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@38647.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@38658.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@38671.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@38706.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@38741.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@38776.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@38811.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@38846.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@38881.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@38916.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@38951.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@38986.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@39021.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@39056.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@39091.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@39126.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@39161.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@39196.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@38646.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@38669.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@38696.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@38731.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@38766.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@38801.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@38836.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@38871.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@38906.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@38941.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@38976.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@39011.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@39046.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@39081.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@39116.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@39151.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@39186.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@39221.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39232.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39233.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39234.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39235.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39236.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39237.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39238.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39239.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39240.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39241.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39242.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39243.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39244.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39245.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39246.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@39263.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@39231.4 FIFOVec.scala 49:42:@39247.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@39282.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@39283.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@39284.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@39285.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@39286.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@39287.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@39288.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@39289.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@39290.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@39291.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@39292.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@39293.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@39294.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@39295.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@39264.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@39298.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@39606.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@39607.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@39608.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@39609.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@39610.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@39611.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@39612.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@39613.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@39614.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@39615.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@39616.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@39617.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@39618.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@39619.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@39620.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@39621.4]
  assign enqCounter_clock = clock; // @[:@38648.4]
  assign enqCounter_reset = reset; // @[:@38649.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@38656.4]
  assign deqCounter_clock = clock; // @[:@38659.4]
  assign deqCounter_reset = reset; // @[:@38660.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@38667.4]
  assign fifos_0_clock = clock; // @[:@38672.4]
  assign fifos_0_reset = reset; // @[:@38673.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@38699.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38701.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38705.4]
  assign fifos_1_clock = clock; // @[:@38707.4]
  assign fifos_1_reset = reset; // @[:@38708.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@38734.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38736.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38740.4]
  assign fifos_2_clock = clock; // @[:@38742.4]
  assign fifos_2_reset = reset; // @[:@38743.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@38769.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38771.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38775.4]
  assign fifos_3_clock = clock; // @[:@38777.4]
  assign fifos_3_reset = reset; // @[:@38778.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@38804.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38806.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38810.4]
  assign fifos_4_clock = clock; // @[:@38812.4]
  assign fifos_4_reset = reset; // @[:@38813.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@38839.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38841.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38845.4]
  assign fifos_5_clock = clock; // @[:@38847.4]
  assign fifos_5_reset = reset; // @[:@38848.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@38874.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38876.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38880.4]
  assign fifos_6_clock = clock; // @[:@38882.4]
  assign fifos_6_reset = reset; // @[:@38883.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@38909.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38911.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38915.4]
  assign fifos_7_clock = clock; // @[:@38917.4]
  assign fifos_7_reset = reset; // @[:@38918.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@38944.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38946.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38950.4]
  assign fifos_8_clock = clock; // @[:@38952.4]
  assign fifos_8_reset = reset; // @[:@38953.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@38979.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38981.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38985.4]
  assign fifos_9_clock = clock; // @[:@38987.4]
  assign fifos_9_reset = reset; // @[:@38988.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@39014.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@39016.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@39020.4]
  assign fifos_10_clock = clock; // @[:@39022.4]
  assign fifos_10_reset = reset; // @[:@39023.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@39049.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@39051.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@39055.4]
  assign fifos_11_clock = clock; // @[:@39057.4]
  assign fifos_11_reset = reset; // @[:@39058.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@39084.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@39086.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@39090.4]
  assign fifos_12_clock = clock; // @[:@39092.4]
  assign fifos_12_reset = reset; // @[:@39093.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@39119.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@39121.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@39125.4]
  assign fifos_13_clock = clock; // @[:@39127.4]
  assign fifos_13_reset = reset; // @[:@39128.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@39154.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@39156.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@39160.4]
  assign fifos_14_clock = clock; // @[:@39162.4]
  assign fifos_14_reset = reset; // @[:@39163.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@39189.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@39191.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@39195.4]
  assign fifos_15_clock = clock; // @[:@39197.4]
  assign fifos_15_reset = reset; // @[:@39198.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@39224.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@39226.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@39230.4]
endmodule
module FFRAM( // @[:@39695.2]
  input        clock, // @[:@39696.4]
  input        reset, // @[:@39697.4]
  input  [1:0] io_raddr, // @[:@39698.4]
  input        io_wen, // @[:@39698.4]
  input  [1:0] io_waddr, // @[:@39698.4]
  input        io_wdata, // @[:@39698.4]
  output       io_rdata, // @[:@39698.4]
  input        io_banks_0_wdata_valid, // @[:@39698.4]
  input        io_banks_0_wdata_bits, // @[:@39698.4]
  input        io_banks_1_wdata_valid, // @[:@39698.4]
  input        io_banks_1_wdata_bits, // @[:@39698.4]
  input        io_banks_2_wdata_valid, // @[:@39698.4]
  input        io_banks_2_wdata_bits, // @[:@39698.4]
  input        io_banks_3_wdata_valid, // @[:@39698.4]
  input        io_banks_3_wdata_bits // @[:@39698.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@39702.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@39703.4]
  wire  _T_89; // @[SRAM.scala 148:25:@39704.4]
  wire  _T_90; // @[SRAM.scala 148:15:@39705.4]
  wire  _T_91; // @[SRAM.scala 149:15:@39707.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@39706.4]
  reg  regs_1; // @[SRAM.scala 145:20:@39713.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@39714.4]
  wire  _T_98; // @[SRAM.scala 148:25:@39715.4]
  wire  _T_99; // @[SRAM.scala 148:15:@39716.4]
  wire  _T_100; // @[SRAM.scala 149:15:@39718.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@39717.4]
  reg  regs_2; // @[SRAM.scala 145:20:@39724.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@39725.4]
  wire  _T_107; // @[SRAM.scala 148:25:@39726.4]
  wire  _T_108; // @[SRAM.scala 148:15:@39727.4]
  wire  _T_109; // @[SRAM.scala 149:15:@39729.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@39728.4]
  reg  regs_3; // @[SRAM.scala 145:20:@39735.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@39736.4]
  wire  _T_116; // @[SRAM.scala 148:25:@39737.4]
  wire  _T_117; // @[SRAM.scala 148:15:@39738.4]
  wire  _T_118; // @[SRAM.scala 149:15:@39740.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@39739.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@39749.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@39749.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@39703.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@39704.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@39705.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@39707.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@39706.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@39714.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@39715.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@39716.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@39718.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@39717.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@39725.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@39726.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@39727.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@39729.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@39728.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@39736.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@39737.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@39738.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@39740.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@39739.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@39749.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@39749.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@39749.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@39751.2]
  input   clock, // @[:@39752.4]
  input   reset, // @[:@39753.4]
  output  io_in_ready, // @[:@39754.4]
  input   io_in_valid, // @[:@39754.4]
  input   io_in_bits, // @[:@39754.4]
  input   io_out_ready, // @[:@39754.4]
  output  io_out_valid, // @[:@39754.4]
  output  io_out_bits // @[:@39754.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@39780.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@39780.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@39780.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@39780.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@39780.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@39780.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@39780.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@39790.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@39790.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@39790.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@39790.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@39790.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@39790.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@39790.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@39805.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@39805.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@39805.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@39805.4]
  wire  writeEn; // @[FIFO.scala 30:29:@39778.4]
  wire  readEn; // @[FIFO.scala 31:29:@39779.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@39800.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@39801.4]
  wire  _T_104; // @[FIFO.scala 45:27:@39802.4]
  wire  empty; // @[FIFO.scala 45:24:@39803.4]
  wire  full; // @[FIFO.scala 46:23:@39804.4]
  wire  _T_157; // @[FIFO.scala 83:17:@39891.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@39892.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@39780.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@39790.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@39805.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@39778.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@39779.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@39801.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@39802.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@39803.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@39804.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@39891.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@39892.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@39898.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@39896.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@39830.4]
  assign enqCounter_clock = clock; // @[:@39781.4]
  assign enqCounter_reset = reset; // @[:@39782.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@39788.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@39789.4]
  assign deqCounter_clock = clock; // @[:@39791.4]
  assign deqCounter_reset = reset; // @[:@39792.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@39798.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@39799.4]
  assign FFRAM_clock = clock; // @[:@39806.4]
  assign FFRAM_reset = reset; // @[:@39807.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@39826.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@39827.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@39828.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@39829.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@39832.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@39831.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@39835.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@39834.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@39838.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@39837.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@39841.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@39840.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@43515.2]
  input   clock, // @[:@43516.4]
  input   reset, // @[:@43517.4]
  output  io_in_ready, // @[:@43518.4]
  input   io_in_valid, // @[:@43518.4]
  input   io_in_bits_0, // @[:@43518.4]
  input   io_out_ready, // @[:@43518.4]
  output  io_out_valid, // @[:@43518.4]
  output  io_out_bits_0, // @[:@43518.4]
  output  io_out_bits_1, // @[:@43518.4]
  output  io_out_bits_2, // @[:@43518.4]
  output  io_out_bits_3, // @[:@43518.4]
  output  io_out_bits_4, // @[:@43518.4]
  output  io_out_bits_5, // @[:@43518.4]
  output  io_out_bits_6, // @[:@43518.4]
  output  io_out_bits_7, // @[:@43518.4]
  output  io_out_bits_8, // @[:@43518.4]
  output  io_out_bits_9, // @[:@43518.4]
  output  io_out_bits_10, // @[:@43518.4]
  output  io_out_bits_11, // @[:@43518.4]
  output  io_out_bits_12, // @[:@43518.4]
  output  io_out_bits_13, // @[:@43518.4]
  output  io_out_bits_14, // @[:@43518.4]
  output  io_out_bits_15 // @[:@43518.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@43522.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@43522.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@43522.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@43522.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@43533.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@43533.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@43533.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@43533.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@43546.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@43581.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@43616.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@43651.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@43686.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@43721.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@43756.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@43791.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@43826.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@43861.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@43896.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@43931.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@43966.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@44001.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@44036.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@44071.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@44071.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@44071.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@44071.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@44071.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@44071.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@44071.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@44071.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@43521.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@43544.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@43571.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@43606.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@43641.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@43676.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@43711.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@43746.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@43781.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@43816.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@43851.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@43886.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@43921.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@43956.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@43991.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@44026.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@44061.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@44096.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44107.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44108.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44109.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44110.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44111.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44112.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44113.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44114.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44115.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44116.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44117.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44118.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44119.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44120.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44121.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@44138.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44122.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@44157.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@44158.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@44159.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@44160.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@44161.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@44162.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@44163.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@44164.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@44165.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@44166.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@44167.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@44168.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@44169.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@44170.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@43522.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@43533.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@43546.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@43581.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@43616.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@43651.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@43686.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@43721.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@43756.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@43791.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@43826.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@43861.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@43896.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@43931.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@43966.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@44001.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@44036.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@44071.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@43521.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@43544.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@43571.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@43606.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@43641.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@43676.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@43711.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@43746.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@43781.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@43816.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@43851.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@43886.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@43921.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@43956.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@43991.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@44026.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@44061.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@44096.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44107.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44108.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44109.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44110.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44111.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44112.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44113.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44114.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44115.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44116.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44117.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44118.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44119.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44120.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44121.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@44138.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@44106.4 FIFOVec.scala 49:42:@44122.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@44157.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@44158.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@44159.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@44160.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@44161.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@44162.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@44163.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@44164.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@44165.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@44166.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@44167.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@44168.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@44169.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@44170.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@44139.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@44173.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@44481.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@44482.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@44483.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@44484.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@44485.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@44486.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@44487.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@44488.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@44489.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@44490.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@44491.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@44492.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@44493.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@44494.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@44495.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@44496.4]
  assign enqCounter_clock = clock; // @[:@43523.4]
  assign enqCounter_reset = reset; // @[:@43524.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@43531.4]
  assign deqCounter_clock = clock; // @[:@43534.4]
  assign deqCounter_reset = reset; // @[:@43535.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@43542.4]
  assign fifos_0_clock = clock; // @[:@43547.4]
  assign fifos_0_reset = reset; // @[:@43548.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@43574.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43576.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43580.4]
  assign fifos_1_clock = clock; // @[:@43582.4]
  assign fifos_1_reset = reset; // @[:@43583.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@43609.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43611.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43615.4]
  assign fifos_2_clock = clock; // @[:@43617.4]
  assign fifos_2_reset = reset; // @[:@43618.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@43644.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43646.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43650.4]
  assign fifos_3_clock = clock; // @[:@43652.4]
  assign fifos_3_reset = reset; // @[:@43653.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@43679.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43681.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43685.4]
  assign fifos_4_clock = clock; // @[:@43687.4]
  assign fifos_4_reset = reset; // @[:@43688.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@43714.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43716.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43720.4]
  assign fifos_5_clock = clock; // @[:@43722.4]
  assign fifos_5_reset = reset; // @[:@43723.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@43749.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43751.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43755.4]
  assign fifos_6_clock = clock; // @[:@43757.4]
  assign fifos_6_reset = reset; // @[:@43758.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@43784.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43786.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43790.4]
  assign fifos_7_clock = clock; // @[:@43792.4]
  assign fifos_7_reset = reset; // @[:@43793.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@43819.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43821.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43825.4]
  assign fifos_8_clock = clock; // @[:@43827.4]
  assign fifos_8_reset = reset; // @[:@43828.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@43854.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43856.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43860.4]
  assign fifos_9_clock = clock; // @[:@43862.4]
  assign fifos_9_reset = reset; // @[:@43863.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@43889.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43891.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43895.4]
  assign fifos_10_clock = clock; // @[:@43897.4]
  assign fifos_10_reset = reset; // @[:@43898.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@43924.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43926.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43930.4]
  assign fifos_11_clock = clock; // @[:@43932.4]
  assign fifos_11_reset = reset; // @[:@43933.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@43959.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43961.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43965.4]
  assign fifos_12_clock = clock; // @[:@43967.4]
  assign fifos_12_reset = reset; // @[:@43968.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@43994.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43996.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44000.4]
  assign fifos_13_clock = clock; // @[:@44002.4]
  assign fifos_13_reset = reset; // @[:@44003.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@44029.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44031.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44035.4]
  assign fifos_14_clock = clock; // @[:@44037.4]
  assign fifos_14_reset = reset; // @[:@44038.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@44064.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44066.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44070.4]
  assign fifos_15_clock = clock; // @[:@44072.4]
  assign fifos_15_reset = reset; // @[:@44073.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@44099.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44101.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44105.4]
endmodule
module FIFOWidthConvert( // @[:@44498.2]
  input         clock, // @[:@44499.4]
  input         reset, // @[:@44500.4]
  output        io_in_ready, // @[:@44501.4]
  input         io_in_valid, // @[:@44501.4]
  input  [31:0] io_in_bits_data_0, // @[:@44501.4]
  input         io_in_bits_strobe, // @[:@44501.4]
  input         io_out_ready, // @[:@44501.4]
  output        io_out_valid, // @[:@44501.4]
  output [31:0] io_out_bits_data_0, // @[:@44501.4]
  output [31:0] io_out_bits_data_1, // @[:@44501.4]
  output [31:0] io_out_bits_data_2, // @[:@44501.4]
  output [31:0] io_out_bits_data_3, // @[:@44501.4]
  output [31:0] io_out_bits_data_4, // @[:@44501.4]
  output [31:0] io_out_bits_data_5, // @[:@44501.4]
  output [31:0] io_out_bits_data_6, // @[:@44501.4]
  output [31:0] io_out_bits_data_7, // @[:@44501.4]
  output [31:0] io_out_bits_data_8, // @[:@44501.4]
  output [31:0] io_out_bits_data_9, // @[:@44501.4]
  output [31:0] io_out_bits_data_10, // @[:@44501.4]
  output [31:0] io_out_bits_data_11, // @[:@44501.4]
  output [31:0] io_out_bits_data_12, // @[:@44501.4]
  output [31:0] io_out_bits_data_13, // @[:@44501.4]
  output [31:0] io_out_bits_data_14, // @[:@44501.4]
  output [31:0] io_out_bits_data_15, // @[:@44501.4]
  output [63:0] io_out_bits_strobe // @[:@44501.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@44503.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@44544.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@44603.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@44609.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@44667.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@44673.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@44674.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@44678.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@44682.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@44686.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@44690.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@44694.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@44698.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@44702.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@44706.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@44710.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@44714.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@44718.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@44722.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@44726.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@44730.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@44734.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@44811.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@44820.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@44829.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@44838.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@44847.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@44856.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@44864.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@44503.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@44544.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@44603.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@44609.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@44667.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@44673.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@44674.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@44678.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@44682.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@44686.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@44690.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@44694.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@44698.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@44702.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@44706.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@44710.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@44714.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@44718.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@44722.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@44726.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@44730.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@44734.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@44811.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@44820.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@44829.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@44838.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@44847.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@44856.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@44864.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@44593.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@44594.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@44643.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@44644.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@44645.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@44646.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@44647.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@44648.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@44649.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@44650.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@44651.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@44652.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@44653.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@44654.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@44655.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@44656.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@44657.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@44658.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@44866.4]
  assign FIFOVec_clock = clock; // @[:@44504.4]
  assign FIFOVec_reset = reset; // @[:@44505.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@44590.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@44589.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@44867.4]
  assign FIFOVec_1_clock = clock; // @[:@44545.4]
  assign FIFOVec_1_reset = reset; // @[:@44546.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@44592.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@44591.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@44868.4]
endmodule
module FFRAM_16( // @[:@44906.2]
  input        clock, // @[:@44907.4]
  input        reset, // @[:@44908.4]
  input  [5:0] io_raddr, // @[:@44909.4]
  input        io_wen, // @[:@44909.4]
  input  [5:0] io_waddr, // @[:@44909.4]
  input        io_wdata, // @[:@44909.4]
  output       io_rdata, // @[:@44909.4]
  input        io_banks_0_wdata_valid, // @[:@44909.4]
  input        io_banks_0_wdata_bits, // @[:@44909.4]
  input        io_banks_1_wdata_valid, // @[:@44909.4]
  input        io_banks_1_wdata_bits, // @[:@44909.4]
  input        io_banks_2_wdata_valid, // @[:@44909.4]
  input        io_banks_2_wdata_bits, // @[:@44909.4]
  input        io_banks_3_wdata_valid, // @[:@44909.4]
  input        io_banks_3_wdata_bits, // @[:@44909.4]
  input        io_banks_4_wdata_valid, // @[:@44909.4]
  input        io_banks_4_wdata_bits, // @[:@44909.4]
  input        io_banks_5_wdata_valid, // @[:@44909.4]
  input        io_banks_5_wdata_bits, // @[:@44909.4]
  input        io_banks_6_wdata_valid, // @[:@44909.4]
  input        io_banks_6_wdata_bits, // @[:@44909.4]
  input        io_banks_7_wdata_valid, // @[:@44909.4]
  input        io_banks_7_wdata_bits, // @[:@44909.4]
  input        io_banks_8_wdata_valid, // @[:@44909.4]
  input        io_banks_8_wdata_bits, // @[:@44909.4]
  input        io_banks_9_wdata_valid, // @[:@44909.4]
  input        io_banks_9_wdata_bits, // @[:@44909.4]
  input        io_banks_10_wdata_valid, // @[:@44909.4]
  input        io_banks_10_wdata_bits, // @[:@44909.4]
  input        io_banks_11_wdata_valid, // @[:@44909.4]
  input        io_banks_11_wdata_bits, // @[:@44909.4]
  input        io_banks_12_wdata_valid, // @[:@44909.4]
  input        io_banks_12_wdata_bits, // @[:@44909.4]
  input        io_banks_13_wdata_valid, // @[:@44909.4]
  input        io_banks_13_wdata_bits, // @[:@44909.4]
  input        io_banks_14_wdata_valid, // @[:@44909.4]
  input        io_banks_14_wdata_bits, // @[:@44909.4]
  input        io_banks_15_wdata_valid, // @[:@44909.4]
  input        io_banks_15_wdata_bits, // @[:@44909.4]
  input        io_banks_16_wdata_valid, // @[:@44909.4]
  input        io_banks_16_wdata_bits, // @[:@44909.4]
  input        io_banks_17_wdata_valid, // @[:@44909.4]
  input        io_banks_17_wdata_bits, // @[:@44909.4]
  input        io_banks_18_wdata_valid, // @[:@44909.4]
  input        io_banks_18_wdata_bits, // @[:@44909.4]
  input        io_banks_19_wdata_valid, // @[:@44909.4]
  input        io_banks_19_wdata_bits, // @[:@44909.4]
  input        io_banks_20_wdata_valid, // @[:@44909.4]
  input        io_banks_20_wdata_bits, // @[:@44909.4]
  input        io_banks_21_wdata_valid, // @[:@44909.4]
  input        io_banks_21_wdata_bits, // @[:@44909.4]
  input        io_banks_22_wdata_valid, // @[:@44909.4]
  input        io_banks_22_wdata_bits, // @[:@44909.4]
  input        io_banks_23_wdata_valid, // @[:@44909.4]
  input        io_banks_23_wdata_bits, // @[:@44909.4]
  input        io_banks_24_wdata_valid, // @[:@44909.4]
  input        io_banks_24_wdata_bits, // @[:@44909.4]
  input        io_banks_25_wdata_valid, // @[:@44909.4]
  input        io_banks_25_wdata_bits, // @[:@44909.4]
  input        io_banks_26_wdata_valid, // @[:@44909.4]
  input        io_banks_26_wdata_bits, // @[:@44909.4]
  input        io_banks_27_wdata_valid, // @[:@44909.4]
  input        io_banks_27_wdata_bits, // @[:@44909.4]
  input        io_banks_28_wdata_valid, // @[:@44909.4]
  input        io_banks_28_wdata_bits, // @[:@44909.4]
  input        io_banks_29_wdata_valid, // @[:@44909.4]
  input        io_banks_29_wdata_bits, // @[:@44909.4]
  input        io_banks_30_wdata_valid, // @[:@44909.4]
  input        io_banks_30_wdata_bits, // @[:@44909.4]
  input        io_banks_31_wdata_valid, // @[:@44909.4]
  input        io_banks_31_wdata_bits, // @[:@44909.4]
  input        io_banks_32_wdata_valid, // @[:@44909.4]
  input        io_banks_32_wdata_bits, // @[:@44909.4]
  input        io_banks_33_wdata_valid, // @[:@44909.4]
  input        io_banks_33_wdata_bits, // @[:@44909.4]
  input        io_banks_34_wdata_valid, // @[:@44909.4]
  input        io_banks_34_wdata_bits, // @[:@44909.4]
  input        io_banks_35_wdata_valid, // @[:@44909.4]
  input        io_banks_35_wdata_bits, // @[:@44909.4]
  input        io_banks_36_wdata_valid, // @[:@44909.4]
  input        io_banks_36_wdata_bits, // @[:@44909.4]
  input        io_banks_37_wdata_valid, // @[:@44909.4]
  input        io_banks_37_wdata_bits, // @[:@44909.4]
  input        io_banks_38_wdata_valid, // @[:@44909.4]
  input        io_banks_38_wdata_bits, // @[:@44909.4]
  input        io_banks_39_wdata_valid, // @[:@44909.4]
  input        io_banks_39_wdata_bits, // @[:@44909.4]
  input        io_banks_40_wdata_valid, // @[:@44909.4]
  input        io_banks_40_wdata_bits, // @[:@44909.4]
  input        io_banks_41_wdata_valid, // @[:@44909.4]
  input        io_banks_41_wdata_bits, // @[:@44909.4]
  input        io_banks_42_wdata_valid, // @[:@44909.4]
  input        io_banks_42_wdata_bits, // @[:@44909.4]
  input        io_banks_43_wdata_valid, // @[:@44909.4]
  input        io_banks_43_wdata_bits, // @[:@44909.4]
  input        io_banks_44_wdata_valid, // @[:@44909.4]
  input        io_banks_44_wdata_bits, // @[:@44909.4]
  input        io_banks_45_wdata_valid, // @[:@44909.4]
  input        io_banks_45_wdata_bits, // @[:@44909.4]
  input        io_banks_46_wdata_valid, // @[:@44909.4]
  input        io_banks_46_wdata_bits, // @[:@44909.4]
  input        io_banks_47_wdata_valid, // @[:@44909.4]
  input        io_banks_47_wdata_bits, // @[:@44909.4]
  input        io_banks_48_wdata_valid, // @[:@44909.4]
  input        io_banks_48_wdata_bits, // @[:@44909.4]
  input        io_banks_49_wdata_valid, // @[:@44909.4]
  input        io_banks_49_wdata_bits, // @[:@44909.4]
  input        io_banks_50_wdata_valid, // @[:@44909.4]
  input        io_banks_50_wdata_bits, // @[:@44909.4]
  input        io_banks_51_wdata_valid, // @[:@44909.4]
  input        io_banks_51_wdata_bits, // @[:@44909.4]
  input        io_banks_52_wdata_valid, // @[:@44909.4]
  input        io_banks_52_wdata_bits, // @[:@44909.4]
  input        io_banks_53_wdata_valid, // @[:@44909.4]
  input        io_banks_53_wdata_bits, // @[:@44909.4]
  input        io_banks_54_wdata_valid, // @[:@44909.4]
  input        io_banks_54_wdata_bits, // @[:@44909.4]
  input        io_banks_55_wdata_valid, // @[:@44909.4]
  input        io_banks_55_wdata_bits, // @[:@44909.4]
  input        io_banks_56_wdata_valid, // @[:@44909.4]
  input        io_banks_56_wdata_bits, // @[:@44909.4]
  input        io_banks_57_wdata_valid, // @[:@44909.4]
  input        io_banks_57_wdata_bits, // @[:@44909.4]
  input        io_banks_58_wdata_valid, // @[:@44909.4]
  input        io_banks_58_wdata_bits, // @[:@44909.4]
  input        io_banks_59_wdata_valid, // @[:@44909.4]
  input        io_banks_59_wdata_bits, // @[:@44909.4]
  input        io_banks_60_wdata_valid, // @[:@44909.4]
  input        io_banks_60_wdata_bits, // @[:@44909.4]
  input        io_banks_61_wdata_valid, // @[:@44909.4]
  input        io_banks_61_wdata_bits, // @[:@44909.4]
  input        io_banks_62_wdata_valid, // @[:@44909.4]
  input        io_banks_62_wdata_bits, // @[:@44909.4]
  input        io_banks_63_wdata_valid, // @[:@44909.4]
  input        io_banks_63_wdata_bits // @[:@44909.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@44913.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@44914.4]
  wire  _T_689; // @[SRAM.scala 148:25:@44915.4]
  wire  _T_690; // @[SRAM.scala 148:15:@44916.4]
  wire  _T_691; // @[SRAM.scala 149:15:@44918.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@44917.4]
  reg  regs_1; // @[SRAM.scala 145:20:@44924.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@44925.4]
  wire  _T_698; // @[SRAM.scala 148:25:@44926.4]
  wire  _T_699; // @[SRAM.scala 148:15:@44927.4]
  wire  _T_700; // @[SRAM.scala 149:15:@44929.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@44928.4]
  reg  regs_2; // @[SRAM.scala 145:20:@44935.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@44936.4]
  wire  _T_707; // @[SRAM.scala 148:25:@44937.4]
  wire  _T_708; // @[SRAM.scala 148:15:@44938.4]
  wire  _T_709; // @[SRAM.scala 149:15:@44940.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@44939.4]
  reg  regs_3; // @[SRAM.scala 145:20:@44946.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@44947.4]
  wire  _T_716; // @[SRAM.scala 148:25:@44948.4]
  wire  _T_717; // @[SRAM.scala 148:15:@44949.4]
  wire  _T_718; // @[SRAM.scala 149:15:@44951.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@44950.4]
  reg  regs_4; // @[SRAM.scala 145:20:@44957.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@44958.4]
  wire  _T_725; // @[SRAM.scala 148:25:@44959.4]
  wire  _T_726; // @[SRAM.scala 148:15:@44960.4]
  wire  _T_727; // @[SRAM.scala 149:15:@44962.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@44961.4]
  reg  regs_5; // @[SRAM.scala 145:20:@44968.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@44969.4]
  wire  _T_734; // @[SRAM.scala 148:25:@44970.4]
  wire  _T_735; // @[SRAM.scala 148:15:@44971.4]
  wire  _T_736; // @[SRAM.scala 149:15:@44973.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@44972.4]
  reg  regs_6; // @[SRAM.scala 145:20:@44979.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@44980.4]
  wire  _T_743; // @[SRAM.scala 148:25:@44981.4]
  wire  _T_744; // @[SRAM.scala 148:15:@44982.4]
  wire  _T_745; // @[SRAM.scala 149:15:@44984.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@44983.4]
  reg  regs_7; // @[SRAM.scala 145:20:@44990.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@44991.4]
  wire  _T_752; // @[SRAM.scala 148:25:@44992.4]
  wire  _T_753; // @[SRAM.scala 148:15:@44993.4]
  wire  _T_754; // @[SRAM.scala 149:15:@44995.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@44994.4]
  reg  regs_8; // @[SRAM.scala 145:20:@45001.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@45002.4]
  wire  _T_761; // @[SRAM.scala 148:25:@45003.4]
  wire  _T_762; // @[SRAM.scala 148:15:@45004.4]
  wire  _T_763; // @[SRAM.scala 149:15:@45006.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@45005.4]
  reg  regs_9; // @[SRAM.scala 145:20:@45012.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@45013.4]
  wire  _T_770; // @[SRAM.scala 148:25:@45014.4]
  wire  _T_771; // @[SRAM.scala 148:15:@45015.4]
  wire  _T_772; // @[SRAM.scala 149:15:@45017.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@45016.4]
  reg  regs_10; // @[SRAM.scala 145:20:@45023.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@45024.4]
  wire  _T_779; // @[SRAM.scala 148:25:@45025.4]
  wire  _T_780; // @[SRAM.scala 148:15:@45026.4]
  wire  _T_781; // @[SRAM.scala 149:15:@45028.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@45027.4]
  reg  regs_11; // @[SRAM.scala 145:20:@45034.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@45035.4]
  wire  _T_788; // @[SRAM.scala 148:25:@45036.4]
  wire  _T_789; // @[SRAM.scala 148:15:@45037.4]
  wire  _T_790; // @[SRAM.scala 149:15:@45039.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@45038.4]
  reg  regs_12; // @[SRAM.scala 145:20:@45045.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@45046.4]
  wire  _T_797; // @[SRAM.scala 148:25:@45047.4]
  wire  _T_798; // @[SRAM.scala 148:15:@45048.4]
  wire  _T_799; // @[SRAM.scala 149:15:@45050.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@45049.4]
  reg  regs_13; // @[SRAM.scala 145:20:@45056.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@45057.4]
  wire  _T_806; // @[SRAM.scala 148:25:@45058.4]
  wire  _T_807; // @[SRAM.scala 148:15:@45059.4]
  wire  _T_808; // @[SRAM.scala 149:15:@45061.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@45060.4]
  reg  regs_14; // @[SRAM.scala 145:20:@45067.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@45068.4]
  wire  _T_815; // @[SRAM.scala 148:25:@45069.4]
  wire  _T_816; // @[SRAM.scala 148:15:@45070.4]
  wire  _T_817; // @[SRAM.scala 149:15:@45072.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@45071.4]
  reg  regs_15; // @[SRAM.scala 145:20:@45078.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@45079.4]
  wire  _T_824; // @[SRAM.scala 148:25:@45080.4]
  wire  _T_825; // @[SRAM.scala 148:15:@45081.4]
  wire  _T_826; // @[SRAM.scala 149:15:@45083.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@45082.4]
  reg  regs_16; // @[SRAM.scala 145:20:@45089.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@45090.4]
  wire  _T_833; // @[SRAM.scala 148:25:@45091.4]
  wire  _T_834; // @[SRAM.scala 148:15:@45092.4]
  wire  _T_835; // @[SRAM.scala 149:15:@45094.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@45093.4]
  reg  regs_17; // @[SRAM.scala 145:20:@45100.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@45101.4]
  wire  _T_842; // @[SRAM.scala 148:25:@45102.4]
  wire  _T_843; // @[SRAM.scala 148:15:@45103.4]
  wire  _T_844; // @[SRAM.scala 149:15:@45105.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@45104.4]
  reg  regs_18; // @[SRAM.scala 145:20:@45111.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@45112.4]
  wire  _T_851; // @[SRAM.scala 148:25:@45113.4]
  wire  _T_852; // @[SRAM.scala 148:15:@45114.4]
  wire  _T_853; // @[SRAM.scala 149:15:@45116.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@45115.4]
  reg  regs_19; // @[SRAM.scala 145:20:@45122.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@45123.4]
  wire  _T_860; // @[SRAM.scala 148:25:@45124.4]
  wire  _T_861; // @[SRAM.scala 148:15:@45125.4]
  wire  _T_862; // @[SRAM.scala 149:15:@45127.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@45126.4]
  reg  regs_20; // @[SRAM.scala 145:20:@45133.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@45134.4]
  wire  _T_869; // @[SRAM.scala 148:25:@45135.4]
  wire  _T_870; // @[SRAM.scala 148:15:@45136.4]
  wire  _T_871; // @[SRAM.scala 149:15:@45138.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@45137.4]
  reg  regs_21; // @[SRAM.scala 145:20:@45144.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@45145.4]
  wire  _T_878; // @[SRAM.scala 148:25:@45146.4]
  wire  _T_879; // @[SRAM.scala 148:15:@45147.4]
  wire  _T_880; // @[SRAM.scala 149:15:@45149.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@45148.4]
  reg  regs_22; // @[SRAM.scala 145:20:@45155.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@45156.4]
  wire  _T_887; // @[SRAM.scala 148:25:@45157.4]
  wire  _T_888; // @[SRAM.scala 148:15:@45158.4]
  wire  _T_889; // @[SRAM.scala 149:15:@45160.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@45159.4]
  reg  regs_23; // @[SRAM.scala 145:20:@45166.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@45167.4]
  wire  _T_896; // @[SRAM.scala 148:25:@45168.4]
  wire  _T_897; // @[SRAM.scala 148:15:@45169.4]
  wire  _T_898; // @[SRAM.scala 149:15:@45171.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@45170.4]
  reg  regs_24; // @[SRAM.scala 145:20:@45177.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@45178.4]
  wire  _T_905; // @[SRAM.scala 148:25:@45179.4]
  wire  _T_906; // @[SRAM.scala 148:15:@45180.4]
  wire  _T_907; // @[SRAM.scala 149:15:@45182.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@45181.4]
  reg  regs_25; // @[SRAM.scala 145:20:@45188.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@45189.4]
  wire  _T_914; // @[SRAM.scala 148:25:@45190.4]
  wire  _T_915; // @[SRAM.scala 148:15:@45191.4]
  wire  _T_916; // @[SRAM.scala 149:15:@45193.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@45192.4]
  reg  regs_26; // @[SRAM.scala 145:20:@45199.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@45200.4]
  wire  _T_923; // @[SRAM.scala 148:25:@45201.4]
  wire  _T_924; // @[SRAM.scala 148:15:@45202.4]
  wire  _T_925; // @[SRAM.scala 149:15:@45204.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@45203.4]
  reg  regs_27; // @[SRAM.scala 145:20:@45210.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@45211.4]
  wire  _T_932; // @[SRAM.scala 148:25:@45212.4]
  wire  _T_933; // @[SRAM.scala 148:15:@45213.4]
  wire  _T_934; // @[SRAM.scala 149:15:@45215.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@45214.4]
  reg  regs_28; // @[SRAM.scala 145:20:@45221.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@45222.4]
  wire  _T_941; // @[SRAM.scala 148:25:@45223.4]
  wire  _T_942; // @[SRAM.scala 148:15:@45224.4]
  wire  _T_943; // @[SRAM.scala 149:15:@45226.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@45225.4]
  reg  regs_29; // @[SRAM.scala 145:20:@45232.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@45233.4]
  wire  _T_950; // @[SRAM.scala 148:25:@45234.4]
  wire  _T_951; // @[SRAM.scala 148:15:@45235.4]
  wire  _T_952; // @[SRAM.scala 149:15:@45237.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@45236.4]
  reg  regs_30; // @[SRAM.scala 145:20:@45243.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@45244.4]
  wire  _T_959; // @[SRAM.scala 148:25:@45245.4]
  wire  _T_960; // @[SRAM.scala 148:15:@45246.4]
  wire  _T_961; // @[SRAM.scala 149:15:@45248.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@45247.4]
  reg  regs_31; // @[SRAM.scala 145:20:@45254.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@45255.4]
  wire  _T_968; // @[SRAM.scala 148:25:@45256.4]
  wire  _T_969; // @[SRAM.scala 148:15:@45257.4]
  wire  _T_970; // @[SRAM.scala 149:15:@45259.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@45258.4]
  reg  regs_32; // @[SRAM.scala 145:20:@45265.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@45266.4]
  wire  _T_977; // @[SRAM.scala 148:25:@45267.4]
  wire  _T_978; // @[SRAM.scala 148:15:@45268.4]
  wire  _T_979; // @[SRAM.scala 149:15:@45270.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@45269.4]
  reg  regs_33; // @[SRAM.scala 145:20:@45276.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@45277.4]
  wire  _T_986; // @[SRAM.scala 148:25:@45278.4]
  wire  _T_987; // @[SRAM.scala 148:15:@45279.4]
  wire  _T_988; // @[SRAM.scala 149:15:@45281.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@45280.4]
  reg  regs_34; // @[SRAM.scala 145:20:@45287.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@45288.4]
  wire  _T_995; // @[SRAM.scala 148:25:@45289.4]
  wire  _T_996; // @[SRAM.scala 148:15:@45290.4]
  wire  _T_997; // @[SRAM.scala 149:15:@45292.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@45291.4]
  reg  regs_35; // @[SRAM.scala 145:20:@45298.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@45299.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@45300.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@45301.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@45303.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@45302.4]
  reg  regs_36; // @[SRAM.scala 145:20:@45309.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@45310.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@45311.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@45312.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@45314.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@45313.4]
  reg  regs_37; // @[SRAM.scala 145:20:@45320.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@45321.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@45322.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@45323.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@45325.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@45324.4]
  reg  regs_38; // @[SRAM.scala 145:20:@45331.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@45332.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@45333.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@45334.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@45336.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@45335.4]
  reg  regs_39; // @[SRAM.scala 145:20:@45342.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@45343.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@45344.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@45345.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@45347.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@45346.4]
  reg  regs_40; // @[SRAM.scala 145:20:@45353.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@45354.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@45355.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@45356.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@45358.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@45357.4]
  reg  regs_41; // @[SRAM.scala 145:20:@45364.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@45365.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@45366.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@45367.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@45369.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@45368.4]
  reg  regs_42; // @[SRAM.scala 145:20:@45375.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@45376.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@45377.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@45378.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@45380.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@45379.4]
  reg  regs_43; // @[SRAM.scala 145:20:@45386.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@45387.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@45388.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@45389.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@45391.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@45390.4]
  reg  regs_44; // @[SRAM.scala 145:20:@45397.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@45398.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@45399.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@45400.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@45402.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@45401.4]
  reg  regs_45; // @[SRAM.scala 145:20:@45408.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@45409.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@45410.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@45411.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@45413.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@45412.4]
  reg  regs_46; // @[SRAM.scala 145:20:@45419.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@45420.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@45421.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@45422.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@45424.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@45423.4]
  reg  regs_47; // @[SRAM.scala 145:20:@45430.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@45431.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@45432.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@45433.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@45435.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@45434.4]
  reg  regs_48; // @[SRAM.scala 145:20:@45441.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@45442.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@45443.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@45444.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@45446.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@45445.4]
  reg  regs_49; // @[SRAM.scala 145:20:@45452.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@45453.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@45454.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@45455.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@45457.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@45456.4]
  reg  regs_50; // @[SRAM.scala 145:20:@45463.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@45464.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@45465.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@45466.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@45468.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@45467.4]
  reg  regs_51; // @[SRAM.scala 145:20:@45474.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@45475.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@45476.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@45477.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@45479.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@45478.4]
  reg  regs_52; // @[SRAM.scala 145:20:@45485.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@45486.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@45487.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@45488.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@45490.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@45489.4]
  reg  regs_53; // @[SRAM.scala 145:20:@45496.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@45497.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@45498.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@45499.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@45501.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@45500.4]
  reg  regs_54; // @[SRAM.scala 145:20:@45507.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@45508.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@45509.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@45510.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@45512.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@45511.4]
  reg  regs_55; // @[SRAM.scala 145:20:@45518.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@45519.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@45520.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@45521.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@45523.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@45522.4]
  reg  regs_56; // @[SRAM.scala 145:20:@45529.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@45530.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@45531.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@45532.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@45534.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@45533.4]
  reg  regs_57; // @[SRAM.scala 145:20:@45540.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@45541.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@45542.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@45543.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@45545.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@45544.4]
  reg  regs_58; // @[SRAM.scala 145:20:@45551.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@45552.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@45553.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@45554.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@45556.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@45555.4]
  reg  regs_59; // @[SRAM.scala 145:20:@45562.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@45563.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@45564.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@45565.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@45567.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@45566.4]
  reg  regs_60; // @[SRAM.scala 145:20:@45573.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@45574.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@45575.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@45576.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@45578.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@45577.4]
  reg  regs_61; // @[SRAM.scala 145:20:@45584.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@45585.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@45586.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@45587.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@45589.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@45588.4]
  reg  regs_62; // @[SRAM.scala 145:20:@45595.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@45596.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@45597.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@45598.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@45600.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@45599.4]
  reg  regs_63; // @[SRAM.scala 145:20:@45606.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@45607.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@45608.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@45609.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@45611.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@45610.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@45680.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@45680.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@44914.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@44915.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@44916.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44918.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@44917.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@44925.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@44926.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@44927.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44929.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@44928.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@44936.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@44937.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@44938.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44940.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@44939.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@44947.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@44948.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@44949.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44951.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@44950.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@44958.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@44959.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@44960.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44962.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@44961.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@44969.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@44970.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@44971.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44973.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@44972.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@44980.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@44981.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@44982.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44984.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@44983.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@44991.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@44992.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@44993.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44995.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@44994.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@45002.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@45003.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@45004.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45006.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@45005.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@45013.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@45014.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@45015.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45017.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@45016.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@45024.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@45025.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@45026.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45028.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@45027.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@45035.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@45036.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@45037.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45039.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@45038.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@45046.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@45047.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@45048.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45050.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@45049.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@45057.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@45058.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@45059.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45061.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@45060.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@45068.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@45069.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@45070.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45072.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@45071.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@45079.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@45080.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@45081.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45083.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@45082.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@45090.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@45091.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@45092.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45094.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@45093.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@45101.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@45102.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@45103.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45105.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@45104.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@45112.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@45113.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@45114.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45116.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@45115.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@45123.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@45124.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@45125.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45127.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@45126.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@45134.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@45135.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@45136.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45138.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@45137.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@45145.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@45146.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@45147.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45149.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@45148.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@45156.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@45157.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@45158.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45160.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@45159.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@45167.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@45168.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@45169.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45171.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@45170.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@45178.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@45179.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@45180.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45182.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@45181.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@45189.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@45190.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@45191.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45193.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@45192.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@45200.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@45201.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@45202.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45204.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@45203.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@45211.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@45212.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@45213.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45215.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@45214.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@45222.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@45223.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@45224.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45226.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@45225.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@45233.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@45234.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@45235.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45237.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@45236.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@45244.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@45245.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@45246.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45248.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@45247.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@45255.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@45256.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@45257.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45259.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@45258.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@45266.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@45267.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@45268.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45270.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@45269.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@45277.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@45278.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@45279.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45281.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@45280.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@45288.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@45289.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@45290.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45292.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@45291.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@45299.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@45300.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@45301.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45303.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@45302.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@45310.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@45311.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@45312.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45314.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@45313.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@45321.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@45322.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@45323.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45325.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@45324.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@45332.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@45333.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@45334.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45336.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@45335.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@45343.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@45344.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@45345.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45347.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@45346.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@45354.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@45355.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@45356.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45358.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@45357.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@45365.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@45366.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@45367.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45369.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@45368.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@45376.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@45377.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@45378.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45380.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@45379.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@45387.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@45388.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@45389.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45391.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@45390.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@45398.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@45399.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@45400.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45402.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@45401.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@45409.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@45410.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@45411.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45413.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@45412.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@45420.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@45421.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@45422.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45424.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@45423.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@45431.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@45432.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@45433.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45435.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@45434.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@45442.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@45443.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@45444.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45446.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@45445.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@45453.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@45454.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@45455.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45457.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@45456.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@45464.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@45465.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@45466.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45468.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@45467.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@45475.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@45476.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@45477.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45479.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@45478.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@45486.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@45487.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@45488.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45490.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@45489.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@45497.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@45498.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@45499.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45501.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@45500.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@45508.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@45509.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@45510.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45512.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@45511.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@45519.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@45520.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@45521.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45523.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@45522.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@45530.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@45531.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@45532.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45534.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@45533.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@45541.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@45542.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@45543.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45545.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@45544.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@45552.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@45553.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@45554.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45556.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@45555.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@45563.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@45564.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@45565.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45567.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@45566.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@45574.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@45575.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@45576.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45578.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@45577.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@45585.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@45586.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@45587.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45589.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@45588.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@45596.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@45597.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@45598.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45600.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@45599.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@45607.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@45608.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@45609.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45611.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@45610.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@45680.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@45680.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@45680.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@45682.2]
  input   clock, // @[:@45683.4]
  input   reset, // @[:@45684.4]
  output  io_in_ready, // @[:@45685.4]
  input   io_in_valid, // @[:@45685.4]
  input   io_in_bits, // @[:@45685.4]
  input   io_out_ready, // @[:@45685.4]
  output  io_out_valid, // @[:@45685.4]
  output  io_out_bits, // @[:@45685.4]
  input   io_banks_0_wdata_valid, // @[:@45685.4]
  input   io_banks_0_wdata_bits, // @[:@45685.4]
  input   io_banks_1_wdata_valid, // @[:@45685.4]
  input   io_banks_1_wdata_bits, // @[:@45685.4]
  input   io_banks_2_wdata_valid, // @[:@45685.4]
  input   io_banks_2_wdata_bits, // @[:@45685.4]
  input   io_banks_3_wdata_valid, // @[:@45685.4]
  input   io_banks_3_wdata_bits, // @[:@45685.4]
  input   io_banks_4_wdata_valid, // @[:@45685.4]
  input   io_banks_4_wdata_bits, // @[:@45685.4]
  input   io_banks_5_wdata_valid, // @[:@45685.4]
  input   io_banks_5_wdata_bits, // @[:@45685.4]
  input   io_banks_6_wdata_valid, // @[:@45685.4]
  input   io_banks_6_wdata_bits, // @[:@45685.4]
  input   io_banks_7_wdata_valid, // @[:@45685.4]
  input   io_banks_7_wdata_bits, // @[:@45685.4]
  input   io_banks_8_wdata_valid, // @[:@45685.4]
  input   io_banks_8_wdata_bits, // @[:@45685.4]
  input   io_banks_9_wdata_valid, // @[:@45685.4]
  input   io_banks_9_wdata_bits, // @[:@45685.4]
  input   io_banks_10_wdata_valid, // @[:@45685.4]
  input   io_banks_10_wdata_bits, // @[:@45685.4]
  input   io_banks_11_wdata_valid, // @[:@45685.4]
  input   io_banks_11_wdata_bits, // @[:@45685.4]
  input   io_banks_12_wdata_valid, // @[:@45685.4]
  input   io_banks_12_wdata_bits, // @[:@45685.4]
  input   io_banks_13_wdata_valid, // @[:@45685.4]
  input   io_banks_13_wdata_bits, // @[:@45685.4]
  input   io_banks_14_wdata_valid, // @[:@45685.4]
  input   io_banks_14_wdata_bits, // @[:@45685.4]
  input   io_banks_15_wdata_valid, // @[:@45685.4]
  input   io_banks_15_wdata_bits, // @[:@45685.4]
  input   io_banks_16_wdata_valid, // @[:@45685.4]
  input   io_banks_16_wdata_bits, // @[:@45685.4]
  input   io_banks_17_wdata_valid, // @[:@45685.4]
  input   io_banks_17_wdata_bits, // @[:@45685.4]
  input   io_banks_18_wdata_valid, // @[:@45685.4]
  input   io_banks_18_wdata_bits, // @[:@45685.4]
  input   io_banks_19_wdata_valid, // @[:@45685.4]
  input   io_banks_19_wdata_bits, // @[:@45685.4]
  input   io_banks_20_wdata_valid, // @[:@45685.4]
  input   io_banks_20_wdata_bits, // @[:@45685.4]
  input   io_banks_21_wdata_valid, // @[:@45685.4]
  input   io_banks_21_wdata_bits, // @[:@45685.4]
  input   io_banks_22_wdata_valid, // @[:@45685.4]
  input   io_banks_22_wdata_bits, // @[:@45685.4]
  input   io_banks_23_wdata_valid, // @[:@45685.4]
  input   io_banks_23_wdata_bits, // @[:@45685.4]
  input   io_banks_24_wdata_valid, // @[:@45685.4]
  input   io_banks_24_wdata_bits, // @[:@45685.4]
  input   io_banks_25_wdata_valid, // @[:@45685.4]
  input   io_banks_25_wdata_bits, // @[:@45685.4]
  input   io_banks_26_wdata_valid, // @[:@45685.4]
  input   io_banks_26_wdata_bits, // @[:@45685.4]
  input   io_banks_27_wdata_valid, // @[:@45685.4]
  input   io_banks_27_wdata_bits, // @[:@45685.4]
  input   io_banks_28_wdata_valid, // @[:@45685.4]
  input   io_banks_28_wdata_bits, // @[:@45685.4]
  input   io_banks_29_wdata_valid, // @[:@45685.4]
  input   io_banks_29_wdata_bits, // @[:@45685.4]
  input   io_banks_30_wdata_valid, // @[:@45685.4]
  input   io_banks_30_wdata_bits, // @[:@45685.4]
  input   io_banks_31_wdata_valid, // @[:@45685.4]
  input   io_banks_31_wdata_bits, // @[:@45685.4]
  input   io_banks_32_wdata_valid, // @[:@45685.4]
  input   io_banks_32_wdata_bits, // @[:@45685.4]
  input   io_banks_33_wdata_valid, // @[:@45685.4]
  input   io_banks_33_wdata_bits, // @[:@45685.4]
  input   io_banks_34_wdata_valid, // @[:@45685.4]
  input   io_banks_34_wdata_bits, // @[:@45685.4]
  input   io_banks_35_wdata_valid, // @[:@45685.4]
  input   io_banks_35_wdata_bits, // @[:@45685.4]
  input   io_banks_36_wdata_valid, // @[:@45685.4]
  input   io_banks_36_wdata_bits, // @[:@45685.4]
  input   io_banks_37_wdata_valid, // @[:@45685.4]
  input   io_banks_37_wdata_bits, // @[:@45685.4]
  input   io_banks_38_wdata_valid, // @[:@45685.4]
  input   io_banks_38_wdata_bits, // @[:@45685.4]
  input   io_banks_39_wdata_valid, // @[:@45685.4]
  input   io_banks_39_wdata_bits, // @[:@45685.4]
  input   io_banks_40_wdata_valid, // @[:@45685.4]
  input   io_banks_40_wdata_bits, // @[:@45685.4]
  input   io_banks_41_wdata_valid, // @[:@45685.4]
  input   io_banks_41_wdata_bits, // @[:@45685.4]
  input   io_banks_42_wdata_valid, // @[:@45685.4]
  input   io_banks_42_wdata_bits, // @[:@45685.4]
  input   io_banks_43_wdata_valid, // @[:@45685.4]
  input   io_banks_43_wdata_bits, // @[:@45685.4]
  input   io_banks_44_wdata_valid, // @[:@45685.4]
  input   io_banks_44_wdata_bits, // @[:@45685.4]
  input   io_banks_45_wdata_valid, // @[:@45685.4]
  input   io_banks_45_wdata_bits, // @[:@45685.4]
  input   io_banks_46_wdata_valid, // @[:@45685.4]
  input   io_banks_46_wdata_bits, // @[:@45685.4]
  input   io_banks_47_wdata_valid, // @[:@45685.4]
  input   io_banks_47_wdata_bits, // @[:@45685.4]
  input   io_banks_48_wdata_valid, // @[:@45685.4]
  input   io_banks_48_wdata_bits, // @[:@45685.4]
  input   io_banks_49_wdata_valid, // @[:@45685.4]
  input   io_banks_49_wdata_bits, // @[:@45685.4]
  input   io_banks_50_wdata_valid, // @[:@45685.4]
  input   io_banks_50_wdata_bits, // @[:@45685.4]
  input   io_banks_51_wdata_valid, // @[:@45685.4]
  input   io_banks_51_wdata_bits, // @[:@45685.4]
  input   io_banks_52_wdata_valid, // @[:@45685.4]
  input   io_banks_52_wdata_bits, // @[:@45685.4]
  input   io_banks_53_wdata_valid, // @[:@45685.4]
  input   io_banks_53_wdata_bits, // @[:@45685.4]
  input   io_banks_54_wdata_valid, // @[:@45685.4]
  input   io_banks_54_wdata_bits, // @[:@45685.4]
  input   io_banks_55_wdata_valid, // @[:@45685.4]
  input   io_banks_55_wdata_bits, // @[:@45685.4]
  input   io_banks_56_wdata_valid, // @[:@45685.4]
  input   io_banks_56_wdata_bits, // @[:@45685.4]
  input   io_banks_57_wdata_valid, // @[:@45685.4]
  input   io_banks_57_wdata_bits, // @[:@45685.4]
  input   io_banks_58_wdata_valid, // @[:@45685.4]
  input   io_banks_58_wdata_bits, // @[:@45685.4]
  input   io_banks_59_wdata_valid, // @[:@45685.4]
  input   io_banks_59_wdata_bits, // @[:@45685.4]
  input   io_banks_60_wdata_valid, // @[:@45685.4]
  input   io_banks_60_wdata_bits, // @[:@45685.4]
  input   io_banks_61_wdata_valid, // @[:@45685.4]
  input   io_banks_61_wdata_bits, // @[:@45685.4]
  input   io_banks_62_wdata_valid, // @[:@45685.4]
  input   io_banks_62_wdata_bits, // @[:@45685.4]
  input   io_banks_63_wdata_valid, // @[:@45685.4]
  input   io_banks_63_wdata_bits // @[:@45685.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@45951.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@45951.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@45951.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@45951.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@45951.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@45961.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@45961.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@45961.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@45961.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@45961.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@45976.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@45976.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@45976.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@45976.4]
  wire  writeEn; // @[FIFO.scala 30:29:@45949.4]
  wire  readEn; // @[FIFO.scala 31:29:@45950.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@45971.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@45972.4]
  wire  _T_824; // @[FIFO.scala 45:27:@45973.4]
  wire  empty; // @[FIFO.scala 45:24:@45974.4]
  wire  full; // @[FIFO.scala 46:23:@45975.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@47142.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@47143.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@45951.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@45961.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@45976.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@45949.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@45950.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@45972.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@45973.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@45974.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@45975.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@47142.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@47143.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@47149.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@47147.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@46181.4]
  assign enqCounter_clock = clock; // @[:@45952.4]
  assign enqCounter_reset = reset; // @[:@45953.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@45959.4]
  assign deqCounter_clock = clock; // @[:@45962.4]
  assign deqCounter_reset = reset; // @[:@45963.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@45969.4]
  assign FFRAM_clock = clock; // @[:@45977.4]
  assign FFRAM_reset = reset; // @[:@45978.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@46177.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@46178.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@46179.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@46180.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@46183.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@46182.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@46186.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@46185.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@46189.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@46188.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@46192.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@46191.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@46195.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@46194.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@46198.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@46197.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@46201.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@46200.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@46204.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@46203.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@46207.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@46206.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@46210.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@46209.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@46213.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@46212.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@46216.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@46215.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@46219.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@46218.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@46222.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@46221.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@46225.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@46224.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@46228.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@46227.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@46231.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@46230.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@46234.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@46233.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@46237.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@46236.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@46240.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@46239.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@46243.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@46242.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@46246.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@46245.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@46249.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@46248.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@46252.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@46251.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@46255.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@46254.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@46258.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@46257.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@46261.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@46260.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@46264.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@46263.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@46267.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@46266.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@46270.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@46269.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@46273.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@46272.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@46276.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@46275.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@46279.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@46278.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@46282.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@46281.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@46285.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@46284.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@46288.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@46287.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@46291.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@46290.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@46294.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@46293.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@46297.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@46296.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@46300.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@46299.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@46303.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@46302.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@46306.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@46305.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@46309.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@46308.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@46312.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@46311.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@46315.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@46314.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@46318.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@46317.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@46321.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@46320.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@46324.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@46323.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@46327.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@46326.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@46330.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@46329.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@46333.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@46332.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@46336.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@46335.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@46339.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@46338.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@46342.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@46341.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@46345.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@46344.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@46348.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@46347.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@46351.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@46350.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@46354.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@46353.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@46357.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@46356.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@46360.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@46359.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@46363.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@46362.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@46366.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@46365.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@46369.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@46368.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@46372.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@46371.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@47151.2]
  input         clock, // @[:@47152.4]
  input         reset, // @[:@47153.4]
  input         io_dram_cmd_ready, // @[:@47154.4]
  output        io_dram_cmd_valid, // @[:@47154.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@47154.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@47154.4]
  input         io_dram_wdata_ready, // @[:@47154.4]
  output        io_dram_wdata_valid, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@47154.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@47154.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@47154.4]
  output        io_dram_wresp_ready, // @[:@47154.4]
  input         io_dram_wresp_valid, // @[:@47154.4]
  output        io_store_cmd_ready, // @[:@47154.4]
  input         io_store_cmd_valid, // @[:@47154.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@47154.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@47154.4]
  output        io_store_data_ready, // @[:@47154.4]
  input         io_store_data_valid, // @[:@47154.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@47154.4]
  input         io_store_data_bits_wstrb, // @[:@47154.4]
  input         io_store_wresp_ready, // @[:@47154.4]
  output        io_store_wresp_valid, // @[:@47154.4]
  output        io_store_wresp_bits // @[:@47154.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@47279.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@47279.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@47279.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@47279.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@47279.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@47279.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@47279.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@47279.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@47279.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@47279.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@47685.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@47685.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@47685.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@47685.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@47685.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@47685.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@47685.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@47685.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@47685.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@47926.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@47926.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@47682.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@47279.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@47685.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@47926.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@47682.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@47679.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@47680.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@47683.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@47715.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@47716.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@47717.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@47718.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@47719.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@47720.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@47721.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@47722.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@47723.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@47724.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@47725.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@47726.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@47727.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@47728.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@47729.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@47730.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@47731.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@47861.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@47862.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@47863.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@47864.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@47865.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@47866.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@47867.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@47868.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@47869.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@47870.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@47871.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@47872.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@47873.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@47874.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@47875.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@47876.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@47877.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@47878.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@47879.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@47880.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@47881.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@47882.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@47883.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@47884.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@47885.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@47886.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@47887.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@47888.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@47889.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@47890.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@47891.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@47892.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@47893.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@47894.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@47895.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@47896.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@47897.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@47898.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@47899.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@47900.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@47901.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@47902.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@47903.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@47904.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@47905.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@47906.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@47907.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@47908.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@47909.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@47910.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@47911.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@47912.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@47913.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@47914.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@47915.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@47916.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@47917.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@47918.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@47919.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@47920.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@47921.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@47922.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@47923.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@47924.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@48193.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@47677.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@47714.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@48194.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@48195.4]
  assign cmd_clock = clock; // @[:@47280.4]
  assign cmd_reset = reset; // @[:@47281.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@47674.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@47676.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@47675.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@47678.4]
  assign wdata_clock = clock; // @[:@47686.4]
  assign wdata_reset = reset; // @[:@47687.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@47711.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@47712.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@47713.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@47925.4]
  assign wresp_clock = clock; // @[:@47927.4]
  assign wresp_reset = reset; // @[:@47928.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@48191.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@48192.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@48196.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@48262.2]
  output        io_in_ready, // @[:@48265.4]
  input         io_in_valid, // @[:@48265.4]
  input  [63:0] io_in_bits_0_addr, // @[:@48265.4]
  input  [31:0] io_in_bits_0_size, // @[:@48265.4]
  input         io_in_bits_0_isWr, // @[:@48265.4]
  input  [31:0] io_in_bits_0_tag, // @[:@48265.4]
  input         io_out_ready, // @[:@48265.4]
  output        io_out_valid, // @[:@48265.4]
  output [63:0] io_out_bits_addr, // @[:@48265.4]
  output [31:0] io_out_bits_size, // @[:@48265.4]
  output        io_out_bits_isWr, // @[:@48265.4]
  output [31:0] io_out_bits_tag // @[:@48265.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@48267.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@48267.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@48276.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@48275.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@48281.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@48280.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@48278.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@48277.4]
endmodule
module MuxPipe_1( // @[:@48283.2]
  output        io_in_ready, // @[:@48286.4]
  input         io_in_valid, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@48286.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@48286.4]
  input         io_in_bits_0_wstrb_0, // @[:@48286.4]
  input         io_in_bits_0_wstrb_1, // @[:@48286.4]
  input         io_in_bits_0_wstrb_2, // @[:@48286.4]
  input         io_in_bits_0_wstrb_3, // @[:@48286.4]
  input         io_in_bits_0_wstrb_4, // @[:@48286.4]
  input         io_in_bits_0_wstrb_5, // @[:@48286.4]
  input         io_in_bits_0_wstrb_6, // @[:@48286.4]
  input         io_in_bits_0_wstrb_7, // @[:@48286.4]
  input         io_in_bits_0_wstrb_8, // @[:@48286.4]
  input         io_in_bits_0_wstrb_9, // @[:@48286.4]
  input         io_in_bits_0_wstrb_10, // @[:@48286.4]
  input         io_in_bits_0_wstrb_11, // @[:@48286.4]
  input         io_in_bits_0_wstrb_12, // @[:@48286.4]
  input         io_in_bits_0_wstrb_13, // @[:@48286.4]
  input         io_in_bits_0_wstrb_14, // @[:@48286.4]
  input         io_in_bits_0_wstrb_15, // @[:@48286.4]
  input         io_in_bits_0_wstrb_16, // @[:@48286.4]
  input         io_in_bits_0_wstrb_17, // @[:@48286.4]
  input         io_in_bits_0_wstrb_18, // @[:@48286.4]
  input         io_in_bits_0_wstrb_19, // @[:@48286.4]
  input         io_in_bits_0_wstrb_20, // @[:@48286.4]
  input         io_in_bits_0_wstrb_21, // @[:@48286.4]
  input         io_in_bits_0_wstrb_22, // @[:@48286.4]
  input         io_in_bits_0_wstrb_23, // @[:@48286.4]
  input         io_in_bits_0_wstrb_24, // @[:@48286.4]
  input         io_in_bits_0_wstrb_25, // @[:@48286.4]
  input         io_in_bits_0_wstrb_26, // @[:@48286.4]
  input         io_in_bits_0_wstrb_27, // @[:@48286.4]
  input         io_in_bits_0_wstrb_28, // @[:@48286.4]
  input         io_in_bits_0_wstrb_29, // @[:@48286.4]
  input         io_in_bits_0_wstrb_30, // @[:@48286.4]
  input         io_in_bits_0_wstrb_31, // @[:@48286.4]
  input         io_in_bits_0_wstrb_32, // @[:@48286.4]
  input         io_in_bits_0_wstrb_33, // @[:@48286.4]
  input         io_in_bits_0_wstrb_34, // @[:@48286.4]
  input         io_in_bits_0_wstrb_35, // @[:@48286.4]
  input         io_in_bits_0_wstrb_36, // @[:@48286.4]
  input         io_in_bits_0_wstrb_37, // @[:@48286.4]
  input         io_in_bits_0_wstrb_38, // @[:@48286.4]
  input         io_in_bits_0_wstrb_39, // @[:@48286.4]
  input         io_in_bits_0_wstrb_40, // @[:@48286.4]
  input         io_in_bits_0_wstrb_41, // @[:@48286.4]
  input         io_in_bits_0_wstrb_42, // @[:@48286.4]
  input         io_in_bits_0_wstrb_43, // @[:@48286.4]
  input         io_in_bits_0_wstrb_44, // @[:@48286.4]
  input         io_in_bits_0_wstrb_45, // @[:@48286.4]
  input         io_in_bits_0_wstrb_46, // @[:@48286.4]
  input         io_in_bits_0_wstrb_47, // @[:@48286.4]
  input         io_in_bits_0_wstrb_48, // @[:@48286.4]
  input         io_in_bits_0_wstrb_49, // @[:@48286.4]
  input         io_in_bits_0_wstrb_50, // @[:@48286.4]
  input         io_in_bits_0_wstrb_51, // @[:@48286.4]
  input         io_in_bits_0_wstrb_52, // @[:@48286.4]
  input         io_in_bits_0_wstrb_53, // @[:@48286.4]
  input         io_in_bits_0_wstrb_54, // @[:@48286.4]
  input         io_in_bits_0_wstrb_55, // @[:@48286.4]
  input         io_in_bits_0_wstrb_56, // @[:@48286.4]
  input         io_in_bits_0_wstrb_57, // @[:@48286.4]
  input         io_in_bits_0_wstrb_58, // @[:@48286.4]
  input         io_in_bits_0_wstrb_59, // @[:@48286.4]
  input         io_in_bits_0_wstrb_60, // @[:@48286.4]
  input         io_in_bits_0_wstrb_61, // @[:@48286.4]
  input         io_in_bits_0_wstrb_62, // @[:@48286.4]
  input         io_in_bits_0_wstrb_63, // @[:@48286.4]
  input         io_out_ready, // @[:@48286.4]
  output        io_out_valid, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_0, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_1, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_2, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_3, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_4, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_5, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_6, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_7, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_8, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_9, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_10, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_11, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_12, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_13, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_14, // @[:@48286.4]
  output [31:0] io_out_bits_wdata_15, // @[:@48286.4]
  output        io_out_bits_wstrb_0, // @[:@48286.4]
  output        io_out_bits_wstrb_1, // @[:@48286.4]
  output        io_out_bits_wstrb_2, // @[:@48286.4]
  output        io_out_bits_wstrb_3, // @[:@48286.4]
  output        io_out_bits_wstrb_4, // @[:@48286.4]
  output        io_out_bits_wstrb_5, // @[:@48286.4]
  output        io_out_bits_wstrb_6, // @[:@48286.4]
  output        io_out_bits_wstrb_7, // @[:@48286.4]
  output        io_out_bits_wstrb_8, // @[:@48286.4]
  output        io_out_bits_wstrb_9, // @[:@48286.4]
  output        io_out_bits_wstrb_10, // @[:@48286.4]
  output        io_out_bits_wstrb_11, // @[:@48286.4]
  output        io_out_bits_wstrb_12, // @[:@48286.4]
  output        io_out_bits_wstrb_13, // @[:@48286.4]
  output        io_out_bits_wstrb_14, // @[:@48286.4]
  output        io_out_bits_wstrb_15, // @[:@48286.4]
  output        io_out_bits_wstrb_16, // @[:@48286.4]
  output        io_out_bits_wstrb_17, // @[:@48286.4]
  output        io_out_bits_wstrb_18, // @[:@48286.4]
  output        io_out_bits_wstrb_19, // @[:@48286.4]
  output        io_out_bits_wstrb_20, // @[:@48286.4]
  output        io_out_bits_wstrb_21, // @[:@48286.4]
  output        io_out_bits_wstrb_22, // @[:@48286.4]
  output        io_out_bits_wstrb_23, // @[:@48286.4]
  output        io_out_bits_wstrb_24, // @[:@48286.4]
  output        io_out_bits_wstrb_25, // @[:@48286.4]
  output        io_out_bits_wstrb_26, // @[:@48286.4]
  output        io_out_bits_wstrb_27, // @[:@48286.4]
  output        io_out_bits_wstrb_28, // @[:@48286.4]
  output        io_out_bits_wstrb_29, // @[:@48286.4]
  output        io_out_bits_wstrb_30, // @[:@48286.4]
  output        io_out_bits_wstrb_31, // @[:@48286.4]
  output        io_out_bits_wstrb_32, // @[:@48286.4]
  output        io_out_bits_wstrb_33, // @[:@48286.4]
  output        io_out_bits_wstrb_34, // @[:@48286.4]
  output        io_out_bits_wstrb_35, // @[:@48286.4]
  output        io_out_bits_wstrb_36, // @[:@48286.4]
  output        io_out_bits_wstrb_37, // @[:@48286.4]
  output        io_out_bits_wstrb_38, // @[:@48286.4]
  output        io_out_bits_wstrb_39, // @[:@48286.4]
  output        io_out_bits_wstrb_40, // @[:@48286.4]
  output        io_out_bits_wstrb_41, // @[:@48286.4]
  output        io_out_bits_wstrb_42, // @[:@48286.4]
  output        io_out_bits_wstrb_43, // @[:@48286.4]
  output        io_out_bits_wstrb_44, // @[:@48286.4]
  output        io_out_bits_wstrb_45, // @[:@48286.4]
  output        io_out_bits_wstrb_46, // @[:@48286.4]
  output        io_out_bits_wstrb_47, // @[:@48286.4]
  output        io_out_bits_wstrb_48, // @[:@48286.4]
  output        io_out_bits_wstrb_49, // @[:@48286.4]
  output        io_out_bits_wstrb_50, // @[:@48286.4]
  output        io_out_bits_wstrb_51, // @[:@48286.4]
  output        io_out_bits_wstrb_52, // @[:@48286.4]
  output        io_out_bits_wstrb_53, // @[:@48286.4]
  output        io_out_bits_wstrb_54, // @[:@48286.4]
  output        io_out_bits_wstrb_55, // @[:@48286.4]
  output        io_out_bits_wstrb_56, // @[:@48286.4]
  output        io_out_bits_wstrb_57, // @[:@48286.4]
  output        io_out_bits_wstrb_58, // @[:@48286.4]
  output        io_out_bits_wstrb_59, // @[:@48286.4]
  output        io_out_bits_wstrb_60, // @[:@48286.4]
  output        io_out_bits_wstrb_61, // @[:@48286.4]
  output        io_out_bits_wstrb_62, // @[:@48286.4]
  output        io_out_bits_wstrb_63 // @[:@48286.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@48288.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@48288.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@48373.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@48372.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@48439.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@48440.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@48441.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@48442.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@48443.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@48444.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@48445.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@48446.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@48447.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@48448.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@48449.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@48450.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@48451.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@48452.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@48453.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@48454.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@48375.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@48376.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@48377.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@48378.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@48379.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@48380.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@48381.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@48382.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@48383.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@48384.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@48385.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@48386.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@48387.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@48388.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@48389.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@48390.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@48391.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@48392.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@48393.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@48394.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@48395.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@48396.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@48397.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@48398.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@48399.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@48400.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@48401.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@48402.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@48403.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@48404.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@48405.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@48406.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@48407.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@48408.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@48409.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@48410.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@48411.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@48412.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@48413.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@48414.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@48415.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@48416.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@48417.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@48418.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@48419.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@48420.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@48421.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@48422.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@48423.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@48424.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@48425.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@48426.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@48427.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@48428.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@48429.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@48430.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@48431.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@48432.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@48433.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@48434.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@48435.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@48436.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@48437.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@48438.4]
endmodule
module ElementCounter( // @[:@48456.2]
  input         clock, // @[:@48457.4]
  input         reset, // @[:@48458.4]
  input         io_reset, // @[:@48459.4]
  input         io_enable, // @[:@48459.4]
  output [31:0] io_out // @[:@48459.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@48461.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@48462.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@48463.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@48468.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@48464.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@48462.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@48463.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@48468.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@48464.4]
  assign io_out = count; // @[Counter.scala 47:10:@48471.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@48473.2]
  input         clock, // @[:@48474.4]
  input         reset, // @[:@48475.4]
  output        io_app_0_cmd_ready, // @[:@48476.4]
  input         io_app_0_cmd_valid, // @[:@48476.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@48476.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@48476.4]
  input         io_app_0_cmd_bits_isWr, // @[:@48476.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@48476.4]
  output        io_app_0_wdata_ready, // @[:@48476.4]
  input         io_app_0_wdata_valid, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@48476.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@48476.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@48476.4]
  input         io_app_0_rresp_ready, // @[:@48476.4]
  input         io_app_0_wresp_ready, // @[:@48476.4]
  output        io_app_0_wresp_valid, // @[:@48476.4]
  input         io_dram_cmd_ready, // @[:@48476.4]
  output        io_dram_cmd_valid, // @[:@48476.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@48476.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@48476.4]
  output        io_dram_cmd_bits_isWr, // @[:@48476.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@48476.4]
  input         io_dram_wdata_ready, // @[:@48476.4]
  output        io_dram_wdata_valid, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@48476.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@48476.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@48476.4]
  output        io_dram_rresp_ready, // @[:@48476.4]
  output        io_dram_wresp_ready, // @[:@48476.4]
  input         io_dram_wresp_valid, // @[:@48476.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@48476.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48705.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48705.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48705.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@48705.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@48705.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48712.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48712.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48712.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48712.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48712.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@48722.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@48722.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@48722.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@48722.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@48722.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@48722.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@48722.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@48722.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@48722.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@48722.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@48722.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@48722.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@48745.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@48745.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@48748.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@48748.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@48748.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@48748.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@48748.4]
  wire  _T_346; // @[package.scala 96:25:@48717.4 package.scala 96:25:@48718.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@48719.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@48721.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@48737.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@48739.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@48742.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@48751.4]
  wire [31:0] _T_365; // @[:@48755.4 :@48756.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@48757.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@48763.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@48766.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@48767.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@48954.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@48961.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@48966.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@48970.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@48971.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@48995.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@48705.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@48712.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@48722.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@48745.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@48748.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@48717.4 package.scala 96:25:@48718.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@48719.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@48721.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@48737.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@48739.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@48742.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@48751.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@48755.4 :@48756.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@48757.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@48763.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@48766.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@48767.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@48954.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@48961.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@48966.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@48970.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@48971.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@48995.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@48968.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@48974.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@48997.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@48857.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@48856.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@48855.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@48853.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@48852.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@48940.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@48924.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@48925.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@48926.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@48927.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@48928.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@48929.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@48930.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@48931.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@48932.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@48933.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@48934.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@48935.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@48936.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@48937.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@48938.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@48939.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@48860.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@48861.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@48862.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@48863.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@48864.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@48865.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@48866.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@48867.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@48868.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@48869.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@48870.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@48871.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@48872.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@48873.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@48874.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@48875.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@48876.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@48877.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@48878.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@48879.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@48880.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@48881.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@48882.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@48883.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@48884.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@48885.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@48886.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@48887.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@48888.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@48889.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@48890.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@48891.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@48892.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@48893.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@48894.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@48895.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@48896.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@48897.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@48898.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@48899.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@48900.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@48901.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@48902.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@48903.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@48904.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@48905.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@48906.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@48907.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@48908.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@48909.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@48910.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@48911.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@48912.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@48913.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@48914.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@48915.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@48916.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@48917.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@48918.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@48919.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@48920.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@48921.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@48922.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@48923.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@49001.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@49004.4]
  assign RetimeWrapper_clock = clock; // @[:@48706.4]
  assign RetimeWrapper_reset = reset; // @[:@48707.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48709.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@48708.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48713.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48714.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48716.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@48715.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@48725.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@48731.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@48730.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@48728.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@48727.4 FringeBundles.scala 115:32:@48744.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@48858.4 StreamArbiter.scala 57:23:@48964.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@48769.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@48836.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@48837.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@48838.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@48839.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@48840.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@48841.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@48842.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@48843.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@48844.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@48845.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@48846.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@48847.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@48848.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@48849.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@48850.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@48851.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@48772.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@48773.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@48774.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@48775.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@48776.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@48777.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@48778.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@48779.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@48780.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@48781.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@48782.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@48783.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@48784.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@48785.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@48786.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@48787.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@48788.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@48789.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@48790.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@48791.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@48792.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@48793.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@48794.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@48795.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@48796.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@48797.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@48798.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@48799.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@48800.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@48801.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@48802.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@48803.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@48804.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@48805.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@48806.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@48807.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@48808.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@48809.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@48810.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@48811.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@48812.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@48813.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@48814.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@48815.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@48816.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@48817.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@48818.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@48819.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@48820.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@48821.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@48822.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@48823.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@48824.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@48825.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@48826.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@48827.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@48828.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@48829.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@48830.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@48831.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@48832.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@48833.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@48834.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@48835.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@48941.4 StreamArbiter.scala 58:25:@48965.4]
  assign elementCtr_clock = clock; // @[:@48749.4]
  assign elementCtr_reset = reset; // @[:@48750.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@48753.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@48752.4]
endmodule
module Counter_72( // @[:@49006.2]
  input         clock, // @[:@49007.4]
  input         reset, // @[:@49008.4]
  input         io_reset, // @[:@49009.4]
  input         io_enable, // @[:@49009.4]
  input  [31:0] io_stride, // @[:@49009.4]
  output [31:0] io_out, // @[:@49009.4]
  output [31:0] io_next // @[:@49009.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@49011.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@49012.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@49013.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@49018.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@49014.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@49012.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@49013.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@49018.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@49014.4]
  assign io_out = count; // @[Counter.scala 25:10:@49021.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@49022.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@49024.2]
  input         clock, // @[:@49025.4]
  input         reset, // @[:@49026.4]
  output        io_in_cmd_ready, // @[:@49027.4]
  input         io_in_cmd_valid, // @[:@49027.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@49027.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@49027.4]
  input         io_in_cmd_bits_isWr, // @[:@49027.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@49027.4]
  output        io_in_wdata_ready, // @[:@49027.4]
  input         io_in_wdata_valid, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@49027.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@49027.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@49027.4]
  input         io_in_rresp_ready, // @[:@49027.4]
  input         io_in_wresp_ready, // @[:@49027.4]
  output        io_in_wresp_valid, // @[:@49027.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@49027.4]
  input         io_out_cmd_ready, // @[:@49027.4]
  output        io_out_cmd_valid, // @[:@49027.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@49027.4]
  output [31:0] io_out_cmd_bits_size, // @[:@49027.4]
  output        io_out_cmd_bits_isWr, // @[:@49027.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@49027.4]
  input         io_out_wdata_ready, // @[:@49027.4]
  output        io_out_wdata_valid, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@49027.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@49027.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@49027.4]
  output        io_out_rresp_ready, // @[:@49027.4]
  output        io_out_wresp_ready, // @[:@49027.4]
  input         io_out_wresp_valid, // @[:@49027.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@49027.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@49141.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@49141.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@49141.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@49141.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@49141.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@49141.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@49141.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@49144.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@49145.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@49146.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@49147.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@49150.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@49150.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@49151.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@49151.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@49152.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@49155.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@49162.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@49166.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@49169.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@49172.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@49183.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@49141.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@49144.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@49145.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@49146.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@49147.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@49150.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@49150.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@49151.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@49151.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@49152.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@49155.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@49162.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@49166.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@49169.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@49172.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@49183.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@49140.4 AXIProtocol.scala 38:19:@49174.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@49133.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@49030.4 AXIProtocol.scala 46:21:@49188.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@49029.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@49139.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@49138.4 AXIProtocol.scala 29:24:@49157.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@49137.4 AXIProtocol.scala 25:24:@49149.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@49135.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@49134.4 FringeBundles.scala 115:32:@49171.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@49132.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@49116.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@49117.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@49118.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@49119.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@49120.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@49121.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@49122.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@49123.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@49124.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@49125.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@49126.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@49127.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@49128.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@49129.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@49130.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@49131.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@49052.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@49053.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@49054.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@49055.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@49056.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@49057.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@49058.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@49059.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@49060.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@49061.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@49062.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@49063.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@49064.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@49065.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@49066.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@49067.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@49068.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@49069.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@49070.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@49071.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@49072.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@49073.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@49074.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@49075.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@49076.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@49077.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@49078.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@49079.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@49080.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@49081.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@49082.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@49083.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@49084.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@49085.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@49086.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@49087.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@49088.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@49089.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@49090.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@49091.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@49092.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@49093.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@49094.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@49095.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@49096.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@49097.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@49098.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@49099.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@49100.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@49101.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@49102.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@49103.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@49104.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@49105.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@49106.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@49107.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@49108.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@49109.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@49110.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@49111.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@49112.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@49113.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@49114.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@49115.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@49050.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@49031.4 AXIProtocol.scala 47:22:@49190.4]
  assign cmdSizeCounter_clock = clock; // @[:@49142.4]
  assign cmdSizeCounter_reset = reset; // @[:@49143.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@49175.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@49176.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@49177.4]
endmodule
module AXICmdIssue( // @[:@49210.2]
  input         clock, // @[:@49211.4]
  input         reset, // @[:@49212.4]
  output        io_in_cmd_ready, // @[:@49213.4]
  input         io_in_cmd_valid, // @[:@49213.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@49213.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@49213.4]
  input         io_in_cmd_bits_isWr, // @[:@49213.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@49213.4]
  output        io_in_wdata_ready, // @[:@49213.4]
  input         io_in_wdata_valid, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@49213.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@49213.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@49213.4]
  input         io_in_rresp_ready, // @[:@49213.4]
  input         io_in_wresp_ready, // @[:@49213.4]
  output        io_in_wresp_valid, // @[:@49213.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@49213.4]
  input         io_out_cmd_ready, // @[:@49213.4]
  output        io_out_cmd_valid, // @[:@49213.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@49213.4]
  output [31:0] io_out_cmd_bits_size, // @[:@49213.4]
  output        io_out_cmd_bits_isWr, // @[:@49213.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@49213.4]
  input         io_out_wdata_ready, // @[:@49213.4]
  output        io_out_wdata_valid, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@49213.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@49213.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@49213.4]
  output        io_out_wdata_bits_wlast, // @[:@49213.4]
  output        io_out_rresp_ready, // @[:@49213.4]
  output        io_out_wresp_ready, // @[:@49213.4]
  input         io_out_wresp_valid, // @[:@49213.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@49213.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@49327.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@49327.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@49327.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@49327.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@49327.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@49327.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@49327.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@49330.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@49331.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@49332.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@49333.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@49334.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@49340.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@49341.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@49336.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@49350.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@49351.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@49327.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@49331.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@49332.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@49333.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@49334.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@49340.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@49341.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@49336.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@49350.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@49351.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@49326.4 AXIProtocol.scala 81:19:@49348.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@49319.4 AXIProtocol.scala 82:21:@49349.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@49216.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@49215.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@49325.4 AXIProtocol.scala 84:20:@49353.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@49324.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@49323.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@49321.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@49320.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@49318.4 AXIProtocol.scala 86:22:@49355.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@49302.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@49303.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@49304.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@49305.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@49306.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@49307.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@49308.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@49309.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@49310.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@49311.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@49312.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@49313.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@49314.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@49315.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@49316.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@49317.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@49238.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@49239.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@49240.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@49241.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@49242.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@49243.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@49244.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@49245.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@49246.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@49247.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@49248.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@49249.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@49250.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@49251.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@49252.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@49253.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@49254.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@49255.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@49256.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@49257.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@49258.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@49259.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@49260.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@49261.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@49262.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@49263.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@49264.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@49265.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@49266.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@49267.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@49268.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@49269.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@49270.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@49271.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@49272.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@49273.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@49274.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@49275.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@49276.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@49277.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@49278.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@49279.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@49280.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@49281.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@49282.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@49283.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@49284.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@49285.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@49286.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@49287.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@49288.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@49289.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@49290.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@49291.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@49292.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@49293.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@49294.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@49295.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@49296.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@49297.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@49298.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@49299.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@49300.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@49301.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@49237.4 AXIProtocol.scala 87:27:@49356.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@49236.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@49217.4]
  assign wdataCounter_clock = clock; // @[:@49328.4]
  assign wdataCounter_reset = reset; // @[:@49329.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@49344.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@49345.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@49346.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@49358.2]
  input         clock, // @[:@49359.4]
  input         reset, // @[:@49360.4]
  input         io_enable, // @[:@49361.4]
  output        io_app_stores_0_cmd_ready, // @[:@49361.4]
  input         io_app_stores_0_cmd_valid, // @[:@49361.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@49361.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@49361.4]
  output        io_app_stores_0_data_ready, // @[:@49361.4]
  input         io_app_stores_0_data_valid, // @[:@49361.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@49361.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@49361.4]
  input         io_app_stores_0_wresp_ready, // @[:@49361.4]
  output        io_app_stores_0_wresp_valid, // @[:@49361.4]
  output        io_app_stores_0_wresp_bits, // @[:@49361.4]
  input         io_dram_cmd_ready, // @[:@49361.4]
  output        io_dram_cmd_valid, // @[:@49361.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@49361.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@49361.4]
  output        io_dram_cmd_bits_isWr, // @[:@49361.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@49361.4]
  input         io_dram_wdata_ready, // @[:@49361.4]
  output        io_dram_wdata_valid, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@49361.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@49361.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@49361.4]
  output        io_dram_wdata_bits_wlast, // @[:@49361.4]
  output        io_dram_rresp_ready, // @[:@49361.4]
  output        io_dram_wresp_ready, // @[:@49361.4]
  input         io_dram_wresp_valid, // @[:@49361.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@49361.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@50247.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@50261.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@50489.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@50604.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@50604.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@50247.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@50261.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@50489.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@50604.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@50260.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@50256.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@50251.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@50250.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@50829.4 DRAMArbiter.scala 100:23:@50832.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@50828.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@50827.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@50825.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@50824.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@50822.4 DRAMArbiter.scala 101:25:@50834.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@50806.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@50807.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@50808.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@50809.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@50810.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@50811.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@50812.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@50813.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@50814.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@50815.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@50816.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@50817.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@50818.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@50819.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@50820.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@50821.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@50742.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@50743.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@50744.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@50745.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@50746.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@50747.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@50748.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@50749.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@50750.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@50751.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@50752.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@50753.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@50754.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@50755.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@50756.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@50757.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@50758.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@50759.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@50760.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@50761.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@50762.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@50763.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@50764.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@50765.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@50766.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@50767.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@50768.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@50769.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@50770.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@50771.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@50772.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@50773.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@50774.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@50775.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@50776.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@50777.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@50778.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@50779.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@50780.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@50781.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@50782.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@50783.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@50784.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@50785.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@50786.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@50787.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@50788.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@50789.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@50790.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@50791.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@50792.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@50793.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@50794.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@50795.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@50796.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@50797.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@50798.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@50799.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@50800.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@50801.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@50802.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@50803.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@50804.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@50805.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@50741.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@50740.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@50721.4]
  assign StreamControllerStore_clock = clock; // @[:@50248.4]
  assign StreamControllerStore_reset = reset; // @[:@50249.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@50376.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@50369.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@50266.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@50259.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@50258.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@50257.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@50255.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@50254.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@50253.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@50252.4]
  assign StreamArbiter_clock = clock; // @[:@50262.4]
  assign StreamArbiter_reset = reset; // @[:@50263.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@50487.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@50486.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@50485.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@50483.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@50482.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@50480.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@50464.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@50465.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@50466.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@50467.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@50468.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@50469.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@50470.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@50471.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@50472.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@50473.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@50474.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@50475.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@50476.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@50477.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@50478.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@50479.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@50400.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@50401.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@50402.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@50403.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@50404.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@50405.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@50406.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@50407.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@50408.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@50409.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@50410.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@50411.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@50412.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@50413.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@50414.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@50415.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@50416.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@50417.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@50418.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@50419.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@50420.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@50421.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@50422.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@50423.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@50424.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@50425.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@50426.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@50427.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@50428.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@50429.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@50430.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@50431.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@50432.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@50433.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@50434.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@50435.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@50436.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@50437.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@50438.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@50439.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@50440.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@50441.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@50442.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@50443.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@50444.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@50445.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@50446.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@50447.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@50448.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@50449.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@50450.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@50451.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@50452.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@50453.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@50454.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@50455.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@50456.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@50457.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@50458.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@50459.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@50460.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@50461.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@50462.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@50463.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@50398.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@50379.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@50603.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@50596.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@50493.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@50492.4]
  assign AXICmdSplit_clock = clock; // @[:@50490.4]
  assign AXICmdSplit_reset = reset; // @[:@50491.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@50602.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@50601.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@50600.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@50598.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@50597.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@50595.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@50579.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@50580.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@50581.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@50582.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@50583.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@50584.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@50585.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@50586.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@50587.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@50588.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@50589.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@50590.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@50591.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@50592.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@50593.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@50594.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@50515.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@50516.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@50517.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@50518.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@50519.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@50520.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@50521.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@50522.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@50523.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@50524.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@50525.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@50526.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@50527.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@50528.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@50529.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@50530.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@50531.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@50532.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@50533.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@50534.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@50535.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@50536.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@50537.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@50538.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@50539.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@50540.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@50541.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@50542.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@50543.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@50544.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@50545.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@50546.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@50547.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@50548.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@50549.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@50550.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@50551.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@50552.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@50553.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@50554.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@50555.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@50556.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@50557.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@50558.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@50559.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@50560.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@50561.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@50562.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@50563.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@50564.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@50565.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@50566.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@50567.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@50568.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@50569.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@50570.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@50571.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@50572.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@50573.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@50574.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@50575.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@50576.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@50577.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@50578.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@50513.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@50494.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@50718.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@50711.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@50608.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@50607.4]
  assign AXICmdIssue_clock = clock; // @[:@50605.4]
  assign AXICmdIssue_reset = reset; // @[:@50606.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@50717.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@50716.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@50715.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@50713.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@50712.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@50710.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@50694.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@50695.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@50696.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@50697.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@50698.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@50699.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@50700.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@50701.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@50702.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@50703.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@50704.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@50705.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@50706.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@50707.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@50708.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@50709.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@50630.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@50631.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@50632.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@50633.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@50634.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@50635.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@50636.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@50637.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@50638.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@50639.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@50640.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@50641.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@50642.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@50643.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@50644.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@50645.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@50646.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@50647.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@50648.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@50649.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@50650.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@50651.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@50652.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@50653.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@50654.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@50655.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@50656.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@50657.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@50658.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@50659.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@50660.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@50661.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@50662.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@50663.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@50664.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@50665.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@50666.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@50667.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@50668.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@50669.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@50670.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@50671.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@50672.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@50673.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@50674.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@50675.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@50676.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@50677.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@50678.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@50679.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@50680.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@50681.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@50682.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@50683.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@50684.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@50685.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@50686.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@50687.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@50688.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@50689.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@50690.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@50691.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@50692.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@50693.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@50628.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@50609.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@50830.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@50823.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@50720.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@50719.4]
endmodule
module DRAMArbiter_1( // @[:@65059.2]
  input         clock, // @[:@65060.4]
  input         reset, // @[:@65061.4]
  input         io_enable, // @[:@65062.4]
  input         io_dram_cmd_ready, // @[:@65062.4]
  output        io_dram_cmd_valid, // @[:@65062.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@65062.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@65062.4]
  output        io_dram_cmd_bits_isWr, // @[:@65062.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@65062.4]
  input         io_dram_wdata_ready, // @[:@65062.4]
  output        io_dram_wdata_valid, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@65062.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@65062.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@65062.4]
  output        io_dram_wdata_bits_wlast, // @[:@65062.4]
  output        io_dram_rresp_ready, // @[:@65062.4]
  output        io_dram_wresp_ready, // @[:@65062.4]
  input         io_dram_wresp_valid, // @[:@65062.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@65062.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@65948.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@65962.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@66190.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@66305.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@66305.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@65948.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@65962.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@66190.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@66305.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@66530.4 DRAMArbiter.scala 100:23:@66533.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@66529.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@66528.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@66526.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@66525.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@66523.4 DRAMArbiter.scala 101:25:@66535.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@66507.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@66508.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@66509.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@66510.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@66511.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@66512.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@66513.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@66514.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@66515.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@66516.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@66517.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@66518.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@66519.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@66520.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@66521.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@66522.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@66443.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@66444.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@66445.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@66446.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@66447.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@66448.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@66449.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@66450.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@66451.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@66452.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@66453.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@66454.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@66455.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@66456.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@66457.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@66458.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@66459.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@66460.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@66461.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@66462.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@66463.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@66464.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@66465.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@66466.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@66467.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@66468.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@66469.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@66470.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@66471.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@66472.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@66473.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@66474.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@66475.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@66476.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@66477.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@66478.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@66479.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@66480.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@66481.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@66482.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@66483.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@66484.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@66485.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@66486.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@66487.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@66488.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@66489.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@66490.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@66491.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@66492.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@66493.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@66494.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@66495.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@66496.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@66497.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@66498.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@66499.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@66500.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@66501.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@66502.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@66503.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@66504.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@66505.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@66506.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@66442.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@66441.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@66422.4]
  assign StreamControllerStore_clock = clock; // @[:@65949.4]
  assign StreamControllerStore_reset = reset; // @[:@65950.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@66077.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@66070.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@65967.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@65960.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@65959.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@65958.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@65956.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@65955.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@65954.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@65953.4]
  assign StreamArbiter_clock = clock; // @[:@65963.4]
  assign StreamArbiter_reset = reset; // @[:@65964.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@66188.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@66187.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@66186.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@66184.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@66183.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@66181.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@66165.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@66166.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@66167.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@66168.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@66169.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@66170.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@66171.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@66172.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@66173.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@66174.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@66175.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@66176.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@66177.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@66178.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@66179.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@66180.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@66101.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@66102.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@66103.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@66104.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@66105.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@66106.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@66107.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@66108.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@66109.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@66110.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@66111.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@66112.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@66113.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@66114.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@66115.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@66116.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@66117.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@66118.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@66119.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@66120.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@66121.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@66122.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@66123.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@66124.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@66125.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@66126.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@66127.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@66128.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@66129.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@66130.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@66131.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@66132.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@66133.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@66134.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@66135.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@66136.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@66137.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@66138.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@66139.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@66140.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@66141.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@66142.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@66143.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@66144.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@66145.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@66146.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@66147.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@66148.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@66149.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@66150.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@66151.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@66152.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@66153.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@66154.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@66155.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@66156.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@66157.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@66158.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@66159.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@66160.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@66161.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@66162.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@66163.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@66164.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@66099.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@66080.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@66304.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@66297.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@66194.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@66193.4]
  assign AXICmdSplit_clock = clock; // @[:@66191.4]
  assign AXICmdSplit_reset = reset; // @[:@66192.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@66303.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@66302.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@66301.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@66299.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@66298.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@66296.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@66280.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@66281.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@66282.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@66283.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@66284.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@66285.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@66286.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@66287.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@66288.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@66289.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@66290.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@66291.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@66292.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@66293.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@66294.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@66295.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@66216.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@66217.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@66218.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@66219.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@66220.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@66221.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@66222.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@66223.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@66224.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@66225.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@66226.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@66227.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@66228.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@66229.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@66230.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@66231.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@66232.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@66233.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@66234.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@66235.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@66236.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@66237.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@66238.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@66239.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@66240.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@66241.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@66242.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@66243.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@66244.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@66245.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@66246.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@66247.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@66248.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@66249.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@66250.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@66251.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@66252.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@66253.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@66254.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@66255.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@66256.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@66257.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@66258.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@66259.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@66260.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@66261.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@66262.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@66263.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@66264.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@66265.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@66266.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@66267.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@66268.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@66269.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@66270.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@66271.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@66272.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@66273.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@66274.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@66275.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@66276.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@66277.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@66278.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@66279.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@66214.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@66195.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@66419.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@66412.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@66309.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@66308.4]
  assign AXICmdIssue_clock = clock; // @[:@66306.4]
  assign AXICmdIssue_reset = reset; // @[:@66307.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@66418.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@66417.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@66416.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@66414.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@66413.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@66411.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@66395.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@66396.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@66397.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@66398.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@66399.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@66400.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@66401.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@66402.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@66403.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@66404.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@66405.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@66406.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@66407.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@66408.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@66409.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@66410.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@66331.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@66332.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@66333.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@66334.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@66335.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@66336.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@66337.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@66338.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@66339.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@66340.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@66341.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@66342.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@66343.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@66344.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@66345.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@66346.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@66347.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@66348.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@66349.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@66350.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@66351.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@66352.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@66353.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@66354.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@66355.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@66356.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@66357.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@66358.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@66359.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@66360.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@66361.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@66362.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@66363.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@66364.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@66365.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@66366.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@66367.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@66368.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@66369.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@66370.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@66371.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@66372.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@66373.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@66374.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@66375.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@66376.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@66377.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@66378.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@66379.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@66380.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@66381.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@66382.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@66383.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@66384.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@66385.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@66386.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@66387.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@66388.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@66389.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@66390.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@66391.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@66392.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@66393.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@66394.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@66329.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@66310.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@66531.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@66524.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@66421.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@66420.4]
endmodule
module DRAMHeap( // @[:@97167.2]
  input         io_accel_0_req_valid, // @[:@97170.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@97170.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@97170.4]
  output        io_accel_0_resp_valid, // @[:@97170.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@97170.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@97170.4]
  output        io_host_0_req_valid, // @[:@97170.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@97170.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@97170.4]
  input         io_host_0_resp_valid, // @[:@97170.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@97170.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@97170.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@97177.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@97179.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@97178.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@97174.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@97173.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@97172.4]
endmodule
module RetimeWrapper_341( // @[:@97193.2]
  input         clock, // @[:@97194.4]
  input         reset, // @[:@97195.4]
  input         io_flow, // @[:@97196.4]
  input  [63:0] io_in, // @[:@97196.4]
  output [63:0] io_out // @[:@97196.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@97198.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@97198.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@97198.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@97198.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@97198.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@97198.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@97198.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@97211.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@97210.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@97209.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@97208.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@97207.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@97205.4]
endmodule
module FringeFF( // @[:@97213.2]
  input         clock, // @[:@97214.4]
  input         reset, // @[:@97215.4]
  input  [63:0] io_in, // @[:@97216.4]
  input         io_reset, // @[:@97216.4]
  output [63:0] io_out, // @[:@97216.4]
  input         io_enable // @[:@97216.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@97219.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@97219.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@97219.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@97219.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@97219.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@97224.4 package.scala 96:25:@97225.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@97230.6]
  RetimeWrapper_341 RetimeWrapper ( // @[package.scala 93:22:@97219.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@97224.4 package.scala 96:25:@97225.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@97230.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@97236.4]
  assign RetimeWrapper_clock = clock; // @[:@97220.4]
  assign RetimeWrapper_reset = reset; // @[:@97221.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@97223.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@97222.4]
endmodule
module MuxN( // @[:@125852.2]
  input  [63:0] io_ins_0, // @[:@125855.4]
  input  [63:0] io_ins_1, // @[:@125855.4]
  input  [63:0] io_ins_2, // @[:@125855.4]
  input  [63:0] io_ins_3, // @[:@125855.4]
  input  [63:0] io_ins_4, // @[:@125855.4]
  input  [63:0] io_ins_5, // @[:@125855.4]
  input  [63:0] io_ins_6, // @[:@125855.4]
  input  [63:0] io_ins_7, // @[:@125855.4]
  input  [63:0] io_ins_8, // @[:@125855.4]
  input  [63:0] io_ins_9, // @[:@125855.4]
  input  [63:0] io_ins_10, // @[:@125855.4]
  input  [63:0] io_ins_11, // @[:@125855.4]
  input  [63:0] io_ins_12, // @[:@125855.4]
  input  [63:0] io_ins_13, // @[:@125855.4]
  input  [63:0] io_ins_14, // @[:@125855.4]
  input  [63:0] io_ins_15, // @[:@125855.4]
  input  [63:0] io_ins_16, // @[:@125855.4]
  input  [63:0] io_ins_17, // @[:@125855.4]
  input  [63:0] io_ins_18, // @[:@125855.4]
  input  [63:0] io_ins_19, // @[:@125855.4]
  input  [63:0] io_ins_20, // @[:@125855.4]
  input  [63:0] io_ins_21, // @[:@125855.4]
  input  [63:0] io_ins_22, // @[:@125855.4]
  input  [63:0] io_ins_23, // @[:@125855.4]
  input  [63:0] io_ins_24, // @[:@125855.4]
  input  [63:0] io_ins_25, // @[:@125855.4]
  input  [63:0] io_ins_26, // @[:@125855.4]
  input  [63:0] io_ins_27, // @[:@125855.4]
  input  [63:0] io_ins_28, // @[:@125855.4]
  input  [63:0] io_ins_29, // @[:@125855.4]
  input  [63:0] io_ins_30, // @[:@125855.4]
  input  [63:0] io_ins_31, // @[:@125855.4]
  input  [63:0] io_ins_32, // @[:@125855.4]
  input  [63:0] io_ins_33, // @[:@125855.4]
  input  [63:0] io_ins_34, // @[:@125855.4]
  input  [63:0] io_ins_35, // @[:@125855.4]
  input  [63:0] io_ins_36, // @[:@125855.4]
  input  [63:0] io_ins_37, // @[:@125855.4]
  input  [63:0] io_ins_38, // @[:@125855.4]
  input  [63:0] io_ins_39, // @[:@125855.4]
  input  [63:0] io_ins_40, // @[:@125855.4]
  input  [63:0] io_ins_41, // @[:@125855.4]
  input  [63:0] io_ins_42, // @[:@125855.4]
  input  [63:0] io_ins_43, // @[:@125855.4]
  input  [63:0] io_ins_44, // @[:@125855.4]
  input  [63:0] io_ins_45, // @[:@125855.4]
  input  [63:0] io_ins_46, // @[:@125855.4]
  input  [63:0] io_ins_47, // @[:@125855.4]
  input  [63:0] io_ins_48, // @[:@125855.4]
  input  [63:0] io_ins_49, // @[:@125855.4]
  input  [63:0] io_ins_50, // @[:@125855.4]
  input  [63:0] io_ins_51, // @[:@125855.4]
  input  [63:0] io_ins_52, // @[:@125855.4]
  input  [63:0] io_ins_53, // @[:@125855.4]
  input  [63:0] io_ins_54, // @[:@125855.4]
  input  [63:0] io_ins_55, // @[:@125855.4]
  input  [63:0] io_ins_56, // @[:@125855.4]
  input  [63:0] io_ins_57, // @[:@125855.4]
  input  [63:0] io_ins_58, // @[:@125855.4]
  input  [63:0] io_ins_59, // @[:@125855.4]
  input  [63:0] io_ins_60, // @[:@125855.4]
  input  [63:0] io_ins_61, // @[:@125855.4]
  input  [63:0] io_ins_62, // @[:@125855.4]
  input  [63:0] io_ins_63, // @[:@125855.4]
  input  [63:0] io_ins_64, // @[:@125855.4]
  input  [63:0] io_ins_65, // @[:@125855.4]
  input  [63:0] io_ins_66, // @[:@125855.4]
  input  [63:0] io_ins_67, // @[:@125855.4]
  input  [63:0] io_ins_68, // @[:@125855.4]
  input  [63:0] io_ins_69, // @[:@125855.4]
  input  [63:0] io_ins_70, // @[:@125855.4]
  input  [63:0] io_ins_71, // @[:@125855.4]
  input  [63:0] io_ins_72, // @[:@125855.4]
  input  [63:0] io_ins_73, // @[:@125855.4]
  input  [63:0] io_ins_74, // @[:@125855.4]
  input  [63:0] io_ins_75, // @[:@125855.4]
  input  [63:0] io_ins_76, // @[:@125855.4]
  input  [63:0] io_ins_77, // @[:@125855.4]
  input  [63:0] io_ins_78, // @[:@125855.4]
  input  [63:0] io_ins_79, // @[:@125855.4]
  input  [63:0] io_ins_80, // @[:@125855.4]
  input  [63:0] io_ins_81, // @[:@125855.4]
  input  [63:0] io_ins_82, // @[:@125855.4]
  input  [63:0] io_ins_83, // @[:@125855.4]
  input  [63:0] io_ins_84, // @[:@125855.4]
  input  [63:0] io_ins_85, // @[:@125855.4]
  input  [63:0] io_ins_86, // @[:@125855.4]
  input  [63:0] io_ins_87, // @[:@125855.4]
  input  [63:0] io_ins_88, // @[:@125855.4]
  input  [63:0] io_ins_89, // @[:@125855.4]
  input  [63:0] io_ins_90, // @[:@125855.4]
  input  [63:0] io_ins_91, // @[:@125855.4]
  input  [63:0] io_ins_92, // @[:@125855.4]
  input  [63:0] io_ins_93, // @[:@125855.4]
  input  [63:0] io_ins_94, // @[:@125855.4]
  input  [63:0] io_ins_95, // @[:@125855.4]
  input  [63:0] io_ins_96, // @[:@125855.4]
  input  [63:0] io_ins_97, // @[:@125855.4]
  input  [63:0] io_ins_98, // @[:@125855.4]
  input  [63:0] io_ins_99, // @[:@125855.4]
  input  [63:0] io_ins_100, // @[:@125855.4]
  input  [63:0] io_ins_101, // @[:@125855.4]
  input  [63:0] io_ins_102, // @[:@125855.4]
  input  [63:0] io_ins_103, // @[:@125855.4]
  input  [63:0] io_ins_104, // @[:@125855.4]
  input  [63:0] io_ins_105, // @[:@125855.4]
  input  [63:0] io_ins_106, // @[:@125855.4]
  input  [63:0] io_ins_107, // @[:@125855.4]
  input  [63:0] io_ins_108, // @[:@125855.4]
  input  [63:0] io_ins_109, // @[:@125855.4]
  input  [63:0] io_ins_110, // @[:@125855.4]
  input  [63:0] io_ins_111, // @[:@125855.4]
  input  [63:0] io_ins_112, // @[:@125855.4]
  input  [63:0] io_ins_113, // @[:@125855.4]
  input  [63:0] io_ins_114, // @[:@125855.4]
  input  [63:0] io_ins_115, // @[:@125855.4]
  input  [63:0] io_ins_116, // @[:@125855.4]
  input  [63:0] io_ins_117, // @[:@125855.4]
  input  [63:0] io_ins_118, // @[:@125855.4]
  input  [63:0] io_ins_119, // @[:@125855.4]
  input  [63:0] io_ins_120, // @[:@125855.4]
  input  [63:0] io_ins_121, // @[:@125855.4]
  input  [63:0] io_ins_122, // @[:@125855.4]
  input  [63:0] io_ins_123, // @[:@125855.4]
  input  [63:0] io_ins_124, // @[:@125855.4]
  input  [63:0] io_ins_125, // @[:@125855.4]
  input  [63:0] io_ins_126, // @[:@125855.4]
  input  [63:0] io_ins_127, // @[:@125855.4]
  input  [63:0] io_ins_128, // @[:@125855.4]
  input  [63:0] io_ins_129, // @[:@125855.4]
  input  [63:0] io_ins_130, // @[:@125855.4]
  input  [63:0] io_ins_131, // @[:@125855.4]
  input  [63:0] io_ins_132, // @[:@125855.4]
  input  [63:0] io_ins_133, // @[:@125855.4]
  input  [63:0] io_ins_134, // @[:@125855.4]
  input  [63:0] io_ins_135, // @[:@125855.4]
  input  [63:0] io_ins_136, // @[:@125855.4]
  input  [63:0] io_ins_137, // @[:@125855.4]
  input  [63:0] io_ins_138, // @[:@125855.4]
  input  [63:0] io_ins_139, // @[:@125855.4]
  input  [63:0] io_ins_140, // @[:@125855.4]
  input  [63:0] io_ins_141, // @[:@125855.4]
  input  [63:0] io_ins_142, // @[:@125855.4]
  input  [63:0] io_ins_143, // @[:@125855.4]
  input  [63:0] io_ins_144, // @[:@125855.4]
  input  [63:0] io_ins_145, // @[:@125855.4]
  input  [63:0] io_ins_146, // @[:@125855.4]
  input  [63:0] io_ins_147, // @[:@125855.4]
  input  [63:0] io_ins_148, // @[:@125855.4]
  input  [63:0] io_ins_149, // @[:@125855.4]
  input  [63:0] io_ins_150, // @[:@125855.4]
  input  [63:0] io_ins_151, // @[:@125855.4]
  input  [63:0] io_ins_152, // @[:@125855.4]
  input  [63:0] io_ins_153, // @[:@125855.4]
  input  [63:0] io_ins_154, // @[:@125855.4]
  input  [63:0] io_ins_155, // @[:@125855.4]
  input  [63:0] io_ins_156, // @[:@125855.4]
  input  [63:0] io_ins_157, // @[:@125855.4]
  input  [63:0] io_ins_158, // @[:@125855.4]
  input  [63:0] io_ins_159, // @[:@125855.4]
  input  [63:0] io_ins_160, // @[:@125855.4]
  input  [63:0] io_ins_161, // @[:@125855.4]
  input  [63:0] io_ins_162, // @[:@125855.4]
  input  [63:0] io_ins_163, // @[:@125855.4]
  input  [63:0] io_ins_164, // @[:@125855.4]
  input  [63:0] io_ins_165, // @[:@125855.4]
  input  [63:0] io_ins_166, // @[:@125855.4]
  input  [63:0] io_ins_167, // @[:@125855.4]
  input  [63:0] io_ins_168, // @[:@125855.4]
  input  [63:0] io_ins_169, // @[:@125855.4]
  input  [63:0] io_ins_170, // @[:@125855.4]
  input  [63:0] io_ins_171, // @[:@125855.4]
  input  [63:0] io_ins_172, // @[:@125855.4]
  input  [63:0] io_ins_173, // @[:@125855.4]
  input  [63:0] io_ins_174, // @[:@125855.4]
  input  [63:0] io_ins_175, // @[:@125855.4]
  input  [63:0] io_ins_176, // @[:@125855.4]
  input  [63:0] io_ins_177, // @[:@125855.4]
  input  [63:0] io_ins_178, // @[:@125855.4]
  input  [63:0] io_ins_179, // @[:@125855.4]
  input  [63:0] io_ins_180, // @[:@125855.4]
  input  [63:0] io_ins_181, // @[:@125855.4]
  input  [63:0] io_ins_182, // @[:@125855.4]
  input  [63:0] io_ins_183, // @[:@125855.4]
  input  [63:0] io_ins_184, // @[:@125855.4]
  input  [63:0] io_ins_185, // @[:@125855.4]
  input  [63:0] io_ins_186, // @[:@125855.4]
  input  [63:0] io_ins_187, // @[:@125855.4]
  input  [63:0] io_ins_188, // @[:@125855.4]
  input  [63:0] io_ins_189, // @[:@125855.4]
  input  [63:0] io_ins_190, // @[:@125855.4]
  input  [63:0] io_ins_191, // @[:@125855.4]
  input  [63:0] io_ins_192, // @[:@125855.4]
  input  [63:0] io_ins_193, // @[:@125855.4]
  input  [63:0] io_ins_194, // @[:@125855.4]
  input  [63:0] io_ins_195, // @[:@125855.4]
  input  [63:0] io_ins_196, // @[:@125855.4]
  input  [63:0] io_ins_197, // @[:@125855.4]
  input  [63:0] io_ins_198, // @[:@125855.4]
  input  [63:0] io_ins_199, // @[:@125855.4]
  input  [63:0] io_ins_200, // @[:@125855.4]
  input  [63:0] io_ins_201, // @[:@125855.4]
  input  [63:0] io_ins_202, // @[:@125855.4]
  input  [63:0] io_ins_203, // @[:@125855.4]
  input  [63:0] io_ins_204, // @[:@125855.4]
  input  [63:0] io_ins_205, // @[:@125855.4]
  input  [63:0] io_ins_206, // @[:@125855.4]
  input  [63:0] io_ins_207, // @[:@125855.4]
  input  [63:0] io_ins_208, // @[:@125855.4]
  input  [63:0] io_ins_209, // @[:@125855.4]
  input  [63:0] io_ins_210, // @[:@125855.4]
  input  [63:0] io_ins_211, // @[:@125855.4]
  input  [63:0] io_ins_212, // @[:@125855.4]
  input  [63:0] io_ins_213, // @[:@125855.4]
  input  [63:0] io_ins_214, // @[:@125855.4]
  input  [63:0] io_ins_215, // @[:@125855.4]
  input  [63:0] io_ins_216, // @[:@125855.4]
  input  [63:0] io_ins_217, // @[:@125855.4]
  input  [63:0] io_ins_218, // @[:@125855.4]
  input  [63:0] io_ins_219, // @[:@125855.4]
  input  [63:0] io_ins_220, // @[:@125855.4]
  input  [63:0] io_ins_221, // @[:@125855.4]
  input  [63:0] io_ins_222, // @[:@125855.4]
  input  [63:0] io_ins_223, // @[:@125855.4]
  input  [63:0] io_ins_224, // @[:@125855.4]
  input  [63:0] io_ins_225, // @[:@125855.4]
  input  [63:0] io_ins_226, // @[:@125855.4]
  input  [63:0] io_ins_227, // @[:@125855.4]
  input  [63:0] io_ins_228, // @[:@125855.4]
  input  [63:0] io_ins_229, // @[:@125855.4]
  input  [63:0] io_ins_230, // @[:@125855.4]
  input  [63:0] io_ins_231, // @[:@125855.4]
  input  [63:0] io_ins_232, // @[:@125855.4]
  input  [63:0] io_ins_233, // @[:@125855.4]
  input  [63:0] io_ins_234, // @[:@125855.4]
  input  [63:0] io_ins_235, // @[:@125855.4]
  input  [63:0] io_ins_236, // @[:@125855.4]
  input  [63:0] io_ins_237, // @[:@125855.4]
  input  [63:0] io_ins_238, // @[:@125855.4]
  input  [63:0] io_ins_239, // @[:@125855.4]
  input  [63:0] io_ins_240, // @[:@125855.4]
  input  [63:0] io_ins_241, // @[:@125855.4]
  input  [63:0] io_ins_242, // @[:@125855.4]
  input  [63:0] io_ins_243, // @[:@125855.4]
  input  [63:0] io_ins_244, // @[:@125855.4]
  input  [63:0] io_ins_245, // @[:@125855.4]
  input  [63:0] io_ins_246, // @[:@125855.4]
  input  [63:0] io_ins_247, // @[:@125855.4]
  input  [63:0] io_ins_248, // @[:@125855.4]
  input  [63:0] io_ins_249, // @[:@125855.4]
  input  [63:0] io_ins_250, // @[:@125855.4]
  input  [63:0] io_ins_251, // @[:@125855.4]
  input  [63:0] io_ins_252, // @[:@125855.4]
  input  [63:0] io_ins_253, // @[:@125855.4]
  input  [63:0] io_ins_254, // @[:@125855.4]
  input  [63:0] io_ins_255, // @[:@125855.4]
  input  [63:0] io_ins_256, // @[:@125855.4]
  input  [63:0] io_ins_257, // @[:@125855.4]
  input  [63:0] io_ins_258, // @[:@125855.4]
  input  [63:0] io_ins_259, // @[:@125855.4]
  input  [63:0] io_ins_260, // @[:@125855.4]
  input  [63:0] io_ins_261, // @[:@125855.4]
  input  [63:0] io_ins_262, // @[:@125855.4]
  input  [63:0] io_ins_263, // @[:@125855.4]
  input  [63:0] io_ins_264, // @[:@125855.4]
  input  [63:0] io_ins_265, // @[:@125855.4]
  input  [63:0] io_ins_266, // @[:@125855.4]
  input  [63:0] io_ins_267, // @[:@125855.4]
  input  [63:0] io_ins_268, // @[:@125855.4]
  input  [63:0] io_ins_269, // @[:@125855.4]
  input  [63:0] io_ins_270, // @[:@125855.4]
  input  [63:0] io_ins_271, // @[:@125855.4]
  input  [63:0] io_ins_272, // @[:@125855.4]
  input  [63:0] io_ins_273, // @[:@125855.4]
  input  [63:0] io_ins_274, // @[:@125855.4]
  input  [63:0] io_ins_275, // @[:@125855.4]
  input  [63:0] io_ins_276, // @[:@125855.4]
  input  [63:0] io_ins_277, // @[:@125855.4]
  input  [63:0] io_ins_278, // @[:@125855.4]
  input  [63:0] io_ins_279, // @[:@125855.4]
  input  [63:0] io_ins_280, // @[:@125855.4]
  input  [63:0] io_ins_281, // @[:@125855.4]
  input  [63:0] io_ins_282, // @[:@125855.4]
  input  [63:0] io_ins_283, // @[:@125855.4]
  input  [63:0] io_ins_284, // @[:@125855.4]
  input  [63:0] io_ins_285, // @[:@125855.4]
  input  [63:0] io_ins_286, // @[:@125855.4]
  input  [63:0] io_ins_287, // @[:@125855.4]
  input  [63:0] io_ins_288, // @[:@125855.4]
  input  [63:0] io_ins_289, // @[:@125855.4]
  input  [63:0] io_ins_290, // @[:@125855.4]
  input  [63:0] io_ins_291, // @[:@125855.4]
  input  [63:0] io_ins_292, // @[:@125855.4]
  input  [63:0] io_ins_293, // @[:@125855.4]
  input  [63:0] io_ins_294, // @[:@125855.4]
  input  [63:0] io_ins_295, // @[:@125855.4]
  input  [63:0] io_ins_296, // @[:@125855.4]
  input  [63:0] io_ins_297, // @[:@125855.4]
  input  [63:0] io_ins_298, // @[:@125855.4]
  input  [63:0] io_ins_299, // @[:@125855.4]
  input  [63:0] io_ins_300, // @[:@125855.4]
  input  [63:0] io_ins_301, // @[:@125855.4]
  input  [63:0] io_ins_302, // @[:@125855.4]
  input  [63:0] io_ins_303, // @[:@125855.4]
  input  [63:0] io_ins_304, // @[:@125855.4]
  input  [63:0] io_ins_305, // @[:@125855.4]
  input  [63:0] io_ins_306, // @[:@125855.4]
  input  [63:0] io_ins_307, // @[:@125855.4]
  input  [63:0] io_ins_308, // @[:@125855.4]
  input  [63:0] io_ins_309, // @[:@125855.4]
  input  [63:0] io_ins_310, // @[:@125855.4]
  input  [63:0] io_ins_311, // @[:@125855.4]
  input  [63:0] io_ins_312, // @[:@125855.4]
  input  [63:0] io_ins_313, // @[:@125855.4]
  input  [63:0] io_ins_314, // @[:@125855.4]
  input  [63:0] io_ins_315, // @[:@125855.4]
  input  [63:0] io_ins_316, // @[:@125855.4]
  input  [63:0] io_ins_317, // @[:@125855.4]
  input  [63:0] io_ins_318, // @[:@125855.4]
  input  [63:0] io_ins_319, // @[:@125855.4]
  input  [63:0] io_ins_320, // @[:@125855.4]
  input  [63:0] io_ins_321, // @[:@125855.4]
  input  [63:0] io_ins_322, // @[:@125855.4]
  input  [63:0] io_ins_323, // @[:@125855.4]
  input  [63:0] io_ins_324, // @[:@125855.4]
  input  [63:0] io_ins_325, // @[:@125855.4]
  input  [63:0] io_ins_326, // @[:@125855.4]
  input  [63:0] io_ins_327, // @[:@125855.4]
  input  [63:0] io_ins_328, // @[:@125855.4]
  input  [63:0] io_ins_329, // @[:@125855.4]
  input  [63:0] io_ins_330, // @[:@125855.4]
  input  [63:0] io_ins_331, // @[:@125855.4]
  input  [63:0] io_ins_332, // @[:@125855.4]
  input  [63:0] io_ins_333, // @[:@125855.4]
  input  [63:0] io_ins_334, // @[:@125855.4]
  input  [63:0] io_ins_335, // @[:@125855.4]
  input  [63:0] io_ins_336, // @[:@125855.4]
  input  [63:0] io_ins_337, // @[:@125855.4]
  input  [63:0] io_ins_338, // @[:@125855.4]
  input  [63:0] io_ins_339, // @[:@125855.4]
  input  [63:0] io_ins_340, // @[:@125855.4]
  input  [63:0] io_ins_341, // @[:@125855.4]
  input  [63:0] io_ins_342, // @[:@125855.4]
  input  [63:0] io_ins_343, // @[:@125855.4]
  input  [63:0] io_ins_344, // @[:@125855.4]
  input  [63:0] io_ins_345, // @[:@125855.4]
  input  [63:0] io_ins_346, // @[:@125855.4]
  input  [63:0] io_ins_347, // @[:@125855.4]
  input  [63:0] io_ins_348, // @[:@125855.4]
  input  [63:0] io_ins_349, // @[:@125855.4]
  input  [63:0] io_ins_350, // @[:@125855.4]
  input  [63:0] io_ins_351, // @[:@125855.4]
  input  [63:0] io_ins_352, // @[:@125855.4]
  input  [63:0] io_ins_353, // @[:@125855.4]
  input  [63:0] io_ins_354, // @[:@125855.4]
  input  [63:0] io_ins_355, // @[:@125855.4]
  input  [63:0] io_ins_356, // @[:@125855.4]
  input  [63:0] io_ins_357, // @[:@125855.4]
  input  [63:0] io_ins_358, // @[:@125855.4]
  input  [63:0] io_ins_359, // @[:@125855.4]
  input  [63:0] io_ins_360, // @[:@125855.4]
  input  [63:0] io_ins_361, // @[:@125855.4]
  input  [63:0] io_ins_362, // @[:@125855.4]
  input  [63:0] io_ins_363, // @[:@125855.4]
  input  [63:0] io_ins_364, // @[:@125855.4]
  input  [63:0] io_ins_365, // @[:@125855.4]
  input  [63:0] io_ins_366, // @[:@125855.4]
  input  [63:0] io_ins_367, // @[:@125855.4]
  input  [63:0] io_ins_368, // @[:@125855.4]
  input  [63:0] io_ins_369, // @[:@125855.4]
  input  [63:0] io_ins_370, // @[:@125855.4]
  input  [63:0] io_ins_371, // @[:@125855.4]
  input  [63:0] io_ins_372, // @[:@125855.4]
  input  [63:0] io_ins_373, // @[:@125855.4]
  input  [63:0] io_ins_374, // @[:@125855.4]
  input  [63:0] io_ins_375, // @[:@125855.4]
  input  [63:0] io_ins_376, // @[:@125855.4]
  input  [63:0] io_ins_377, // @[:@125855.4]
  input  [63:0] io_ins_378, // @[:@125855.4]
  input  [63:0] io_ins_379, // @[:@125855.4]
  input  [63:0] io_ins_380, // @[:@125855.4]
  input  [63:0] io_ins_381, // @[:@125855.4]
  input  [63:0] io_ins_382, // @[:@125855.4]
  input  [63:0] io_ins_383, // @[:@125855.4]
  input  [63:0] io_ins_384, // @[:@125855.4]
  input  [63:0] io_ins_385, // @[:@125855.4]
  input  [63:0] io_ins_386, // @[:@125855.4]
  input  [63:0] io_ins_387, // @[:@125855.4]
  input  [63:0] io_ins_388, // @[:@125855.4]
  input  [63:0] io_ins_389, // @[:@125855.4]
  input  [63:0] io_ins_390, // @[:@125855.4]
  input  [63:0] io_ins_391, // @[:@125855.4]
  input  [63:0] io_ins_392, // @[:@125855.4]
  input  [63:0] io_ins_393, // @[:@125855.4]
  input  [63:0] io_ins_394, // @[:@125855.4]
  input  [63:0] io_ins_395, // @[:@125855.4]
  input  [63:0] io_ins_396, // @[:@125855.4]
  input  [63:0] io_ins_397, // @[:@125855.4]
  input  [63:0] io_ins_398, // @[:@125855.4]
  input  [63:0] io_ins_399, // @[:@125855.4]
  input  [63:0] io_ins_400, // @[:@125855.4]
  input  [63:0] io_ins_401, // @[:@125855.4]
  input  [63:0] io_ins_402, // @[:@125855.4]
  input  [63:0] io_ins_403, // @[:@125855.4]
  input  [63:0] io_ins_404, // @[:@125855.4]
  input  [63:0] io_ins_405, // @[:@125855.4]
  input  [63:0] io_ins_406, // @[:@125855.4]
  input  [63:0] io_ins_407, // @[:@125855.4]
  input  [63:0] io_ins_408, // @[:@125855.4]
  input  [63:0] io_ins_409, // @[:@125855.4]
  input  [63:0] io_ins_410, // @[:@125855.4]
  input  [63:0] io_ins_411, // @[:@125855.4]
  input  [63:0] io_ins_412, // @[:@125855.4]
  input  [63:0] io_ins_413, // @[:@125855.4]
  input  [63:0] io_ins_414, // @[:@125855.4]
  input  [63:0] io_ins_415, // @[:@125855.4]
  input  [63:0] io_ins_416, // @[:@125855.4]
  input  [63:0] io_ins_417, // @[:@125855.4]
  input  [63:0] io_ins_418, // @[:@125855.4]
  input  [63:0] io_ins_419, // @[:@125855.4]
  input  [63:0] io_ins_420, // @[:@125855.4]
  input  [63:0] io_ins_421, // @[:@125855.4]
  input  [63:0] io_ins_422, // @[:@125855.4]
  input  [63:0] io_ins_423, // @[:@125855.4]
  input  [63:0] io_ins_424, // @[:@125855.4]
  input  [63:0] io_ins_425, // @[:@125855.4]
  input  [63:0] io_ins_426, // @[:@125855.4]
  input  [63:0] io_ins_427, // @[:@125855.4]
  input  [63:0] io_ins_428, // @[:@125855.4]
  input  [63:0] io_ins_429, // @[:@125855.4]
  input  [63:0] io_ins_430, // @[:@125855.4]
  input  [63:0] io_ins_431, // @[:@125855.4]
  input  [63:0] io_ins_432, // @[:@125855.4]
  input  [63:0] io_ins_433, // @[:@125855.4]
  input  [63:0] io_ins_434, // @[:@125855.4]
  input  [63:0] io_ins_435, // @[:@125855.4]
  input  [63:0] io_ins_436, // @[:@125855.4]
  input  [63:0] io_ins_437, // @[:@125855.4]
  input  [63:0] io_ins_438, // @[:@125855.4]
  input  [63:0] io_ins_439, // @[:@125855.4]
  input  [63:0] io_ins_440, // @[:@125855.4]
  input  [63:0] io_ins_441, // @[:@125855.4]
  input  [63:0] io_ins_442, // @[:@125855.4]
  input  [63:0] io_ins_443, // @[:@125855.4]
  input  [63:0] io_ins_444, // @[:@125855.4]
  input  [63:0] io_ins_445, // @[:@125855.4]
  input  [63:0] io_ins_446, // @[:@125855.4]
  input  [63:0] io_ins_447, // @[:@125855.4]
  input  [63:0] io_ins_448, // @[:@125855.4]
  input  [63:0] io_ins_449, // @[:@125855.4]
  input  [63:0] io_ins_450, // @[:@125855.4]
  input  [63:0] io_ins_451, // @[:@125855.4]
  input  [63:0] io_ins_452, // @[:@125855.4]
  input  [63:0] io_ins_453, // @[:@125855.4]
  input  [63:0] io_ins_454, // @[:@125855.4]
  input  [63:0] io_ins_455, // @[:@125855.4]
  input  [63:0] io_ins_456, // @[:@125855.4]
  input  [63:0] io_ins_457, // @[:@125855.4]
  input  [63:0] io_ins_458, // @[:@125855.4]
  input  [63:0] io_ins_459, // @[:@125855.4]
  input  [63:0] io_ins_460, // @[:@125855.4]
  input  [63:0] io_ins_461, // @[:@125855.4]
  input  [63:0] io_ins_462, // @[:@125855.4]
  input  [63:0] io_ins_463, // @[:@125855.4]
  input  [63:0] io_ins_464, // @[:@125855.4]
  input  [63:0] io_ins_465, // @[:@125855.4]
  input  [63:0] io_ins_466, // @[:@125855.4]
  input  [63:0] io_ins_467, // @[:@125855.4]
  input  [63:0] io_ins_468, // @[:@125855.4]
  input  [63:0] io_ins_469, // @[:@125855.4]
  input  [63:0] io_ins_470, // @[:@125855.4]
  input  [63:0] io_ins_471, // @[:@125855.4]
  input  [63:0] io_ins_472, // @[:@125855.4]
  input  [63:0] io_ins_473, // @[:@125855.4]
  input  [63:0] io_ins_474, // @[:@125855.4]
  input  [63:0] io_ins_475, // @[:@125855.4]
  input  [63:0] io_ins_476, // @[:@125855.4]
  input  [63:0] io_ins_477, // @[:@125855.4]
  input  [63:0] io_ins_478, // @[:@125855.4]
  input  [63:0] io_ins_479, // @[:@125855.4]
  input  [63:0] io_ins_480, // @[:@125855.4]
  input  [63:0] io_ins_481, // @[:@125855.4]
  input  [63:0] io_ins_482, // @[:@125855.4]
  input  [63:0] io_ins_483, // @[:@125855.4]
  input  [63:0] io_ins_484, // @[:@125855.4]
  input  [63:0] io_ins_485, // @[:@125855.4]
  input  [63:0] io_ins_486, // @[:@125855.4]
  input  [63:0] io_ins_487, // @[:@125855.4]
  input  [63:0] io_ins_488, // @[:@125855.4]
  input  [63:0] io_ins_489, // @[:@125855.4]
  input  [63:0] io_ins_490, // @[:@125855.4]
  input  [63:0] io_ins_491, // @[:@125855.4]
  input  [63:0] io_ins_492, // @[:@125855.4]
  input  [63:0] io_ins_493, // @[:@125855.4]
  input  [63:0] io_ins_494, // @[:@125855.4]
  input  [63:0] io_ins_495, // @[:@125855.4]
  input  [63:0] io_ins_496, // @[:@125855.4]
  input  [63:0] io_ins_497, // @[:@125855.4]
  input  [63:0] io_ins_498, // @[:@125855.4]
  input  [63:0] io_ins_499, // @[:@125855.4]
  input  [63:0] io_ins_500, // @[:@125855.4]
  input  [63:0] io_ins_501, // @[:@125855.4]
  input  [63:0] io_ins_502, // @[:@125855.4]
  input  [8:0]  io_sel, // @[:@125855.4]
  output [63:0] io_out // @[:@125855.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@125857.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@125857.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@125857.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@125857.4]
endmodule
module RegFile( // @[:@125859.2]
  input         clock, // @[:@125860.4]
  input         reset, // @[:@125861.4]
  input  [31:0] io_raddr, // @[:@125862.4]
  input         io_wen, // @[:@125862.4]
  input  [31:0] io_waddr, // @[:@125862.4]
  input  [63:0] io_wdata, // @[:@125862.4]
  output [63:0] io_rdata, // @[:@125862.4]
  input         io_reset, // @[:@125862.4]
  output [63:0] io_argIns_0, // @[:@125862.4]
  output [63:0] io_argIns_1, // @[:@125862.4]
  output [63:0] io_argIns_2, // @[:@125862.4]
  output [63:0] io_argIns_3, // @[:@125862.4]
  input         io_argOuts_0_valid, // @[:@125862.4]
  input  [63:0] io_argOuts_0_bits, // @[:@125862.4]
  input         io_argOuts_1_valid, // @[:@125862.4]
  input  [63:0] io_argOuts_1_bits // @[:@125862.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@127872.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@127872.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@127872.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@127872.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@127872.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@127872.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@127884.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@127884.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@127884.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@127884.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@127884.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@127884.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@127903.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@127903.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@127903.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@127903.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@127903.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@127903.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@127915.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@127915.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@127915.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@127915.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@127915.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@127915.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@127927.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@127927.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@127927.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@127927.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@127927.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@127927.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@127941.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@127941.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@127941.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@127941.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@127941.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@127941.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@127955.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@127955.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@127955.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@127955.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@127955.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@127955.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@127969.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@127969.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@127969.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@127969.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@127969.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@127969.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@127983.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@127983.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@127983.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@127983.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@127983.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@127983.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@127997.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@127997.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@127997.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@127997.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@127997.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@127997.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@128011.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@128011.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@128011.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@128011.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@128011.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@128011.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@128025.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@128025.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@128025.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@128025.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@128025.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@128025.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@128039.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@128039.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@128039.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@128039.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@128039.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@128039.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@128053.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@128053.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@128053.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@128053.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@128053.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@128053.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@128067.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@128067.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@128067.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@128067.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@128067.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@128067.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@128081.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@128081.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@128081.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@128081.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@128081.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@128081.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@128095.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@128095.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@128095.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@128095.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@128095.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@128095.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@128109.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@128109.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@128109.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@128109.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@128109.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@128109.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@128123.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@128123.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@128123.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@128123.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@128123.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@128123.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@128137.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@128137.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@128137.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@128137.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@128137.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@128137.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@128151.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@128151.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@128151.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@128151.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@128151.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@128151.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@128165.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@128165.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@128165.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@128165.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@128165.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@128165.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@128179.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@128179.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@128179.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@128179.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@128179.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@128179.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@128193.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@128193.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@128193.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@128193.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@128193.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@128193.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@128207.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@128207.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@128207.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@128207.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@128207.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@128207.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@128221.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@128221.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@128221.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@128221.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@128221.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@128221.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@128235.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@128235.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@128235.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@128235.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@128235.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@128235.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@128249.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@128249.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@128249.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@128249.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@128249.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@128249.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@128263.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@128263.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@128263.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@128263.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@128263.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@128263.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@128277.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@128277.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@128277.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@128277.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@128277.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@128277.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@128291.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@128291.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@128291.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@128291.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@128291.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@128291.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@128305.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@128305.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@128305.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@128305.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@128305.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@128305.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@128319.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@128319.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@128319.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@128319.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@128319.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@128319.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@128333.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@128333.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@128333.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@128333.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@128333.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@128333.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@128347.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@128347.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@128347.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@128347.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@128347.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@128347.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@128361.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@128361.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@128361.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@128361.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@128361.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@128361.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@128375.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@128375.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@128375.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@128375.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@128375.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@128375.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@128389.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@128389.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@128389.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@128389.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@128389.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@128389.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@128403.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@128403.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@128403.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@128403.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@128403.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@128403.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@128417.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@128417.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@128417.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@128417.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@128417.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@128417.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@128431.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@128431.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@128431.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@128431.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@128431.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@128431.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@128445.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@128445.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@128445.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@128445.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@128445.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@128445.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@128459.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@128459.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@128459.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@128459.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@128459.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@128459.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@128473.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@128473.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@128473.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@128473.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@128473.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@128473.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@128487.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@128487.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@128487.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@128487.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@128487.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@128487.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@128501.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@128501.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@128501.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@128501.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@128501.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@128501.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@128515.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@128515.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@128515.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@128515.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@128515.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@128515.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@128529.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@128529.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@128529.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@128529.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@128529.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@128529.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@128543.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@128543.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@128543.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@128543.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@128543.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@128543.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@128557.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@128557.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@128557.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@128557.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@128557.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@128557.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@128571.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@128571.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@128571.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@128571.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@128571.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@128571.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@128585.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@128585.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@128585.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@128585.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@128585.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@128585.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@128599.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@128599.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@128599.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@128599.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@128599.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@128599.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@128613.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@128613.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@128613.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@128613.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@128613.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@128613.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@128627.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@128627.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@128627.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@128627.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@128627.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@128627.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@128641.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@128641.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@128641.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@128641.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@128641.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@128641.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@128655.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@128655.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@128655.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@128655.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@128655.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@128655.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@128669.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@128669.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@128669.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@128669.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@128669.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@128669.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@128683.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@128683.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@128683.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@128683.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@128683.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@128683.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@128697.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@128697.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@128697.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@128697.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@128697.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@128697.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@128711.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@128711.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@128711.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@128711.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@128711.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@128711.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@128725.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@128725.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@128725.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@128725.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@128725.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@128725.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@128739.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@128739.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@128739.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@128739.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@128739.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@128739.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@128753.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@128753.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@128753.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@128753.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@128753.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@128753.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@128767.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@128767.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@128767.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@128767.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@128767.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@128767.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@128781.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@128781.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@128781.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@128781.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@128781.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@128781.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@128795.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@128795.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@128795.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@128795.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@128795.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@128795.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@128809.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@128809.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@128809.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@128809.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@128809.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@128809.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@128823.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@128823.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@128823.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@128823.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@128823.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@128823.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@128837.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@128837.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@128837.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@128837.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@128837.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@128837.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@128851.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@128851.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@128851.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@128851.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@128851.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@128851.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@128865.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@128865.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@128865.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@128865.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@128865.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@128865.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@128879.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@128879.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@128879.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@128879.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@128879.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@128879.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@128893.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@128893.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@128893.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@128893.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@128893.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@128893.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@128907.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@128907.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@128907.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@128907.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@128907.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@128907.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@128921.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@128921.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@128921.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@128921.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@128921.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@128921.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@128935.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@128935.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@128935.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@128935.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@128935.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@128935.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@128949.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@128949.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@128949.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@128949.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@128949.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@128949.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@128963.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@128963.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@128963.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@128963.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@128963.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@128963.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@128977.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@128977.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@128977.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@128977.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@128977.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@128977.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@128991.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@128991.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@128991.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@128991.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@128991.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@128991.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@129005.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@129005.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@129005.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@129005.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@129005.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@129005.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@129019.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@129019.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@129019.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@129019.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@129019.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@129019.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@129033.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@129033.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@129033.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@129033.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@129033.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@129033.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@129047.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@129047.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@129047.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@129047.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@129047.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@129047.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@129061.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@129061.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@129061.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@129061.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@129061.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@129061.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@129075.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@129075.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@129075.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@129075.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@129075.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@129075.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@129089.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@129089.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@129089.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@129089.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@129089.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@129089.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@129103.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@129103.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@129103.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@129103.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@129103.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@129103.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@129117.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@129117.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@129117.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@129117.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@129117.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@129117.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@129131.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@129131.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@129131.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@129131.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@129131.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@129131.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@129145.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@129145.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@129145.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@129145.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@129145.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@129145.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@129159.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@129159.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@129159.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@129159.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@129159.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@129159.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@129173.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@129173.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@129173.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@129173.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@129173.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@129173.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@129187.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@129187.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@129187.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@129187.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@129187.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@129187.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@129201.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@129201.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@129201.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@129201.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@129201.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@129201.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@129215.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@129215.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@129215.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@129215.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@129215.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@129215.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@129229.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@129229.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@129229.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@129229.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@129229.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@129229.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@129243.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@129243.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@129243.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@129243.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@129243.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@129243.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@129257.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@129257.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@129257.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@129257.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@129257.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@129257.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@129271.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@129271.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@129271.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@129271.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@129271.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@129271.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@129285.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@129285.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@129285.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@129285.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@129285.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@129285.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@129299.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@129299.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@129299.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@129299.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@129299.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@129299.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@129313.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@129313.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@129313.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@129313.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@129313.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@129313.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@129327.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@129327.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@129327.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@129327.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@129327.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@129327.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@129341.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@129341.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@129341.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@129341.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@129341.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@129341.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@129355.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@129355.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@129355.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@129355.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@129355.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@129355.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@129369.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@129369.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@129369.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@129369.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@129369.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@129369.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@129383.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@129383.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@129383.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@129383.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@129383.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@129383.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@129397.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@129397.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@129397.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@129397.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@129397.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@129397.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@129411.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@129411.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@129411.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@129411.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@129411.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@129411.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@129425.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@129425.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@129425.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@129425.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@129425.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@129425.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@129439.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@129439.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@129439.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@129439.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@129439.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@129439.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@129453.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@129453.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@129453.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@129453.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@129453.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@129453.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@129467.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@129467.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@129467.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@129467.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@129467.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@129467.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@129481.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@129481.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@129481.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@129481.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@129481.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@129481.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@129495.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@129495.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@129495.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@129495.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@129495.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@129495.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@129509.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@129509.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@129509.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@129509.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@129509.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@129509.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@129523.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@129523.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@129523.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@129523.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@129523.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@129523.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@129537.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@129537.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@129537.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@129537.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@129537.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@129537.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@129551.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@129551.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@129551.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@129551.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@129551.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@129551.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@129565.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@129565.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@129565.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@129565.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@129565.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@129565.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@129579.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@129579.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@129579.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@129579.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@129579.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@129579.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@129593.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@129593.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@129593.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@129593.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@129593.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@129593.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@129607.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@129607.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@129607.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@129607.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@129607.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@129607.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@129621.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@129621.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@129621.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@129621.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@129621.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@129621.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@129635.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@129635.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@129635.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@129635.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@129635.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@129635.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@129649.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@129649.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@129649.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@129649.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@129649.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@129649.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@129663.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@129663.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@129663.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@129663.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@129663.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@129663.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@129677.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@129677.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@129677.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@129677.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@129677.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@129677.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@129691.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@129691.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@129691.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@129691.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@129691.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@129691.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@129705.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@129705.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@129705.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@129705.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@129705.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@129705.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@129719.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@129719.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@129719.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@129719.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@129719.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@129719.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@129733.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@129733.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@129733.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@129733.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@129733.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@129733.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@129747.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@129747.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@129747.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@129747.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@129747.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@129747.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@129761.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@129761.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@129761.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@129761.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@129761.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@129761.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@129775.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@129775.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@129775.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@129775.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@129775.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@129775.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@129789.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@129789.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@129789.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@129789.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@129789.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@129789.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@129803.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@129803.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@129803.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@129803.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@129803.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@129803.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@129817.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@129817.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@129817.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@129817.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@129817.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@129817.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@129831.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@129831.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@129831.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@129831.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@129831.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@129831.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@129845.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@129845.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@129845.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@129845.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@129845.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@129845.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@129859.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@129859.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@129859.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@129859.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@129859.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@129859.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@129873.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@129873.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@129873.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@129873.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@129873.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@129873.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@129887.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@129887.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@129887.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@129887.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@129887.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@129887.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@129901.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@129901.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@129901.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@129901.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@129901.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@129901.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@129915.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@129915.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@129915.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@129915.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@129915.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@129915.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@129929.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@129929.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@129929.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@129929.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@129929.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@129929.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@129943.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@129943.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@129943.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@129943.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@129943.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@129943.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@129957.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@129957.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@129957.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@129957.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@129957.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@129957.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@129971.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@129971.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@129971.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@129971.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@129971.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@129971.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@129985.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@129985.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@129985.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@129985.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@129985.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@129985.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@129999.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@129999.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@129999.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@129999.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@129999.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@129999.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@130013.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@130013.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@130013.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@130013.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@130013.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@130013.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@130027.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@130027.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@130027.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@130027.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@130027.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@130027.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@130041.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@130041.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@130041.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@130041.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@130041.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@130041.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@130055.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@130055.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@130055.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@130055.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@130055.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@130055.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@130069.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@130069.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@130069.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@130069.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@130069.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@130069.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@130083.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@130083.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@130083.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@130083.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@130083.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@130083.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@130097.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@130097.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@130097.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@130097.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@130097.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@130097.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@130111.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@130111.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@130111.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@130111.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@130111.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@130111.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@130125.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@130125.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@130125.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@130125.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@130125.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@130125.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@130139.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@130139.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@130139.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@130139.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@130139.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@130139.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@130153.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@130153.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@130153.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@130153.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@130153.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@130153.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@130167.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@130167.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@130167.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@130167.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@130167.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@130167.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@130181.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@130181.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@130181.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@130181.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@130181.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@130181.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@130195.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@130195.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@130195.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@130195.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@130195.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@130195.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@130209.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@130209.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@130209.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@130209.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@130209.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@130209.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@130223.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@130223.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@130223.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@130223.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@130223.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@130223.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@130237.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@130237.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@130237.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@130237.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@130237.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@130237.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@130251.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@130251.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@130251.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@130251.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@130251.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@130251.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@130265.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@130265.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@130265.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@130265.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@130265.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@130265.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@130279.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@130279.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@130279.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@130279.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@130279.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@130279.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@130293.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@130293.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@130293.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@130293.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@130293.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@130293.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@130307.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@130307.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@130307.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@130307.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@130307.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@130307.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@130321.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@130321.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@130321.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@130321.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@130321.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@130321.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@130335.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@130335.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@130335.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@130335.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@130335.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@130335.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@130349.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@130349.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@130349.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@130349.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@130349.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@130349.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@130363.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@130363.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@130363.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@130363.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@130363.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@130363.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@130377.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@130377.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@130377.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@130377.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@130377.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@130377.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@130391.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@130391.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@130391.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@130391.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@130391.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@130391.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@130405.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@130405.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@130405.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@130405.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@130405.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@130405.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@130419.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@130419.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@130419.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@130419.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@130419.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@130419.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@130433.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@130433.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@130433.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@130433.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@130433.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@130433.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@130447.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@130447.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@130447.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@130447.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@130447.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@130447.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@130461.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@130461.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@130461.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@130461.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@130461.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@130461.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@130475.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@130475.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@130475.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@130475.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@130475.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@130475.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@130489.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@130489.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@130489.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@130489.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@130489.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@130489.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@130503.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@130503.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@130503.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@130503.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@130503.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@130503.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@130517.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@130517.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@130517.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@130517.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@130517.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@130517.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@130531.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@130531.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@130531.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@130531.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@130531.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@130531.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@130545.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@130545.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@130545.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@130545.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@130545.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@130545.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@130559.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@130559.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@130559.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@130559.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@130559.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@130559.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@130573.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@130573.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@130573.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@130573.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@130573.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@130573.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@130587.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@130587.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@130587.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@130587.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@130587.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@130587.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@130601.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@130601.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@130601.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@130601.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@130601.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@130601.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@130615.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@130615.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@130615.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@130615.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@130615.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@130615.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@130629.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@130629.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@130629.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@130629.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@130629.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@130629.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@130643.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@130643.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@130643.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@130643.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@130643.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@130643.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@130657.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@130657.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@130657.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@130657.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@130657.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@130657.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@130671.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@130671.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@130671.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@130671.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@130671.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@130671.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@130685.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@130685.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@130685.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@130685.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@130685.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@130685.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@130699.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@130699.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@130699.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@130699.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@130699.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@130699.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@130713.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@130713.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@130713.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@130713.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@130713.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@130713.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@130727.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@130727.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@130727.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@130727.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@130727.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@130727.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@130741.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@130741.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@130741.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@130741.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@130741.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@130741.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@130755.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@130755.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@130755.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@130755.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@130755.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@130755.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@130769.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@130769.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@130769.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@130769.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@130769.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@130769.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@130783.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@130783.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@130783.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@130783.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@130783.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@130783.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@130797.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@130797.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@130797.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@130797.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@130797.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@130797.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@130811.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@130811.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@130811.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@130811.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@130811.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@130811.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@130825.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@130825.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@130825.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@130825.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@130825.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@130825.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@130839.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@130839.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@130839.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@130839.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@130839.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@130839.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@130853.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@130853.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@130853.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@130853.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@130853.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@130853.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@130867.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@130867.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@130867.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@130867.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@130867.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@130867.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@130881.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@130881.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@130881.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@130881.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@130881.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@130881.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@130895.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@130895.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@130895.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@130895.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@130895.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@130895.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@130909.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@130909.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@130909.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@130909.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@130909.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@130909.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@130923.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@130923.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@130923.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@130923.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@130923.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@130923.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@130937.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@130937.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@130937.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@130937.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@130937.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@130937.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@130951.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@130951.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@130951.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@130951.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@130951.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@130951.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@130965.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@130965.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@130965.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@130965.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@130965.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@130965.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@130979.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@130979.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@130979.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@130979.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@130979.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@130979.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@130993.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@130993.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@130993.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@130993.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@130993.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@130993.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@131007.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@131007.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@131007.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@131007.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@131007.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@131007.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@131021.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@131021.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@131021.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@131021.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@131021.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@131021.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@131035.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@131035.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@131035.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@131035.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@131035.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@131035.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@131049.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@131049.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@131049.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@131049.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@131049.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@131049.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@131063.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@131063.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@131063.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@131063.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@131063.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@131063.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@131077.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@131077.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@131077.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@131077.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@131077.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@131077.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@131091.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@131091.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@131091.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@131091.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@131091.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@131091.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@131105.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@131105.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@131105.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@131105.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@131105.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@131105.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@131119.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@131119.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@131119.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@131119.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@131119.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@131119.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@131133.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@131133.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@131133.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@131133.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@131133.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@131133.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@131147.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@131147.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@131147.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@131147.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@131147.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@131147.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@131161.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@131161.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@131161.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@131161.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@131161.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@131161.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@131175.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@131175.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@131175.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@131175.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@131175.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@131175.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@131189.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@131189.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@131189.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@131189.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@131189.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@131189.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@131203.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@131203.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@131203.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@131203.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@131203.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@131203.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@131217.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@131217.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@131217.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@131217.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@131217.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@131217.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@131231.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@131231.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@131231.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@131231.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@131231.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@131231.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@131245.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@131245.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@131245.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@131245.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@131245.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@131245.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@131259.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@131259.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@131259.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@131259.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@131259.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@131259.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@131273.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@131273.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@131273.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@131273.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@131273.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@131273.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@131287.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@131287.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@131287.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@131287.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@131287.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@131287.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@131301.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@131301.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@131301.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@131301.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@131301.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@131301.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@131315.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@131315.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@131315.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@131315.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@131315.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@131315.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@131329.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@131329.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@131329.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@131329.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@131329.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@131329.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@131343.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@131343.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@131343.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@131343.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@131343.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@131343.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@131357.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@131357.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@131357.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@131357.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@131357.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@131357.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@131371.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@131371.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@131371.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@131371.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@131371.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@131371.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@131385.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@131385.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@131385.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@131385.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@131385.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@131385.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@131399.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@131399.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@131399.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@131399.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@131399.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@131399.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@131413.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@131413.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@131413.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@131413.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@131413.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@131413.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@131427.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@131427.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@131427.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@131427.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@131427.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@131427.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@131441.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@131441.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@131441.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@131441.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@131441.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@131441.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@131455.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@131455.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@131455.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@131455.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@131455.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@131455.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@131469.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@131469.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@131469.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@131469.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@131469.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@131469.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@131483.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@131483.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@131483.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@131483.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@131483.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@131483.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@131497.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@131497.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@131497.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@131497.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@131497.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@131497.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@131511.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@131511.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@131511.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@131511.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@131511.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@131511.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@131525.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@131525.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@131525.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@131525.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@131525.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@131525.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@131539.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@131539.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@131539.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@131539.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@131539.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@131539.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@131553.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@131553.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@131553.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@131553.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@131553.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@131553.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@131567.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@131567.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@131567.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@131567.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@131567.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@131567.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@131581.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@131581.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@131581.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@131581.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@131581.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@131581.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@131595.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@131595.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@131595.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@131595.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@131595.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@131595.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@131609.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@131609.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@131609.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@131609.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@131609.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@131609.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@131623.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@131623.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@131623.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@131623.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@131623.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@131623.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@131637.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@131637.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@131637.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@131637.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@131637.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@131637.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@131651.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@131651.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@131651.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@131651.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@131651.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@131651.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@131665.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@131665.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@131665.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@131665.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@131665.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@131665.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@131679.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@131679.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@131679.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@131679.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@131679.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@131679.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@131693.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@131693.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@131693.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@131693.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@131693.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@131693.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@131707.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@131707.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@131707.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@131707.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@131707.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@131707.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@131721.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@131721.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@131721.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@131721.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@131721.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@131721.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@131735.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@131735.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@131735.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@131735.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@131735.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@131735.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@131749.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@131749.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@131749.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@131749.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@131749.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@131749.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@131763.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@131763.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@131763.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@131763.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@131763.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@131763.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@131777.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@131777.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@131777.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@131777.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@131777.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@131777.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@131791.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@131791.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@131791.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@131791.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@131791.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@131791.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@131805.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@131805.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@131805.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@131805.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@131805.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@131805.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@131819.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@131819.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@131819.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@131819.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@131819.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@131819.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@131833.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@131833.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@131833.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@131833.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@131833.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@131833.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@131847.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@131847.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@131847.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@131847.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@131847.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@131847.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@131861.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@131861.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@131861.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@131861.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@131861.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@131861.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@131875.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@131875.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@131875.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@131875.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@131875.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@131875.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@131889.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@131889.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@131889.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@131889.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@131889.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@131889.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@131903.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@131903.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@131903.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@131903.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@131903.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@131903.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@131917.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@131917.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@131917.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@131917.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@131917.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@131917.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@131931.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@131931.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@131931.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@131931.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@131931.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@131931.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@131945.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@131945.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@131945.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@131945.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@131945.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@131945.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@131959.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@131959.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@131959.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@131959.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@131959.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@131959.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@131973.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@131973.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@131973.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@131973.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@131973.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@131973.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@131987.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@131987.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@131987.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@131987.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@131987.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@131987.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@132001.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@132001.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@132001.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@132001.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@132001.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@132001.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@132015.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@132015.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@132015.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@132015.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@132015.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@132015.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@132029.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@132029.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@132029.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@132029.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@132029.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@132029.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@132043.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@132043.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@132043.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@132043.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@132043.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@132043.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@132057.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@132057.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@132057.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@132057.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@132057.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@132057.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@132071.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@132071.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@132071.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@132071.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@132071.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@132071.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@132085.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@132085.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@132085.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@132085.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@132085.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@132085.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@132099.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@132099.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@132099.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@132099.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@132099.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@132099.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@132113.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@132113.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@132113.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@132113.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@132113.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@132113.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@132127.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@132127.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@132127.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@132127.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@132127.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@132127.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@132141.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@132141.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@132141.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@132141.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@132141.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@132141.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@132155.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@132155.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@132155.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@132155.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@132155.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@132155.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@132169.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@132169.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@132169.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@132169.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@132169.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@132169.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@132183.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@132183.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@132183.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@132183.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@132183.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@132183.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@132197.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@132197.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@132197.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@132197.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@132197.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@132197.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@132211.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@132211.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@132211.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@132211.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@132211.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@132211.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@132225.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@132225.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@132225.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@132225.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@132225.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@132225.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@132239.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@132239.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@132239.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@132239.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@132239.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@132239.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@132253.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@132253.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@132253.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@132253.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@132253.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@132253.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@132267.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@132267.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@132267.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@132267.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@132267.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@132267.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@132281.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@132281.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@132281.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@132281.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@132281.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@132281.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@132295.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@132295.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@132295.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@132295.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@132295.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@132295.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@132309.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@132309.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@132309.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@132309.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@132309.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@132309.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@132323.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@132323.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@132323.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@132323.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@132323.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@132323.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@132337.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@132337.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@132337.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@132337.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@132337.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@132337.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@132351.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@132351.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@132351.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@132351.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@132351.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@132351.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@132365.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@132365.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@132365.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@132365.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@132365.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@132365.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@132379.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@132379.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@132379.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@132379.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@132379.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@132379.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@132393.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@132393.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@132393.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@132393.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@132393.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@132393.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@132407.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@132407.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@132407.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@132407.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@132407.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@132407.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@132421.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@132421.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@132421.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@132421.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@132421.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@132421.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@132435.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@132435.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@132435.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@132435.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@132435.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@132435.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@132449.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@132449.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@132449.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@132449.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@132449.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@132449.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@132463.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@132463.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@132463.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@132463.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@132463.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@132463.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@132477.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@132477.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@132477.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@132477.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@132477.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@132477.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@132491.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@132491.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@132491.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@132491.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@132491.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@132491.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@132505.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@132505.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@132505.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@132505.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@132505.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@132505.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@132519.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@132519.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@132519.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@132519.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@132519.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@132519.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@132533.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@132533.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@132533.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@132533.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@132533.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@132533.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@132547.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@132547.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@132547.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@132547.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@132547.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@132547.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@132561.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@132561.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@132561.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@132561.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@132561.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@132561.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@132575.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@132575.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@132575.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@132575.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@132575.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@132575.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@132589.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@132589.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@132589.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@132589.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@132589.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@132589.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@132603.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@132603.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@132603.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@132603.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@132603.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@132603.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@132617.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@132617.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@132617.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@132617.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@132617.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@132617.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@132631.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@132631.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@132631.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@132631.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@132631.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@132631.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@132645.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@132645.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@132645.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@132645.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@132645.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@132645.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@132659.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@132659.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@132659.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@132659.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@132659.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@132659.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@132673.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@132673.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@132673.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@132673.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@132673.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@132673.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@132687.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@132687.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@132687.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@132687.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@132687.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@132687.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@132701.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@132701.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@132701.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@132701.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@132701.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@132701.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@132715.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@132715.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@132715.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@132715.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@132715.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@132715.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@132729.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@132729.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@132729.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@132729.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@132729.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@132729.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@132743.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@132743.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@132743.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@132743.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@132743.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@132743.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@132757.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@132757.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@132757.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@132757.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@132757.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@132757.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@132771.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@132771.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@132771.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@132771.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@132771.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@132771.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@132785.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@132785.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@132785.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@132785.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@132785.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@132785.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@132799.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@132799.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@132799.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@132799.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@132799.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@132799.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@132813.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@132813.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@132813.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@132813.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@132813.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@132813.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@132827.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@132827.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@132827.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@132827.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@132827.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@132827.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@132841.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@132841.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@132841.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@132841.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@132841.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@132841.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@132855.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@132855.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@132855.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@132855.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@132855.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@132855.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@132869.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@132869.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@132869.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@132869.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@132869.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@132869.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@132883.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@132883.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@132883.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@132883.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@132883.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@132883.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@132897.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@132897.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@132897.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@132897.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@132897.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@132897.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@132911.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@132911.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@132911.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@132911.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@132911.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@132911.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@132925.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@132925.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@132925.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@132925.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@132925.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@132925.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@132939.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@132939.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@132939.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@132939.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@132939.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@132939.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@132953.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@132953.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@132953.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@132953.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@132953.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@132953.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@132967.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@132967.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@132967.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@132967.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@132967.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@132967.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@132981.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@132981.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@132981.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@132981.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@132981.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@132981.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@132995.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@132995.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@132995.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@132995.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@132995.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@132995.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@133009.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@133009.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@133009.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@133009.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@133009.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@133009.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@133023.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@133023.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@133023.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@133023.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@133023.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@133023.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@133037.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@133037.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@133037.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@133037.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@133037.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@133037.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@133051.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@133051.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@133051.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@133051.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@133051.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@133051.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@133065.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@133065.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@133065.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@133065.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@133065.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@133065.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@133079.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@133079.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@133079.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@133079.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@133079.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@133079.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@133093.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@133093.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@133093.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@133093.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@133093.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@133093.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@133107.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@133107.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@133107.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@133107.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@133107.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@133107.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@133121.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@133121.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@133121.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@133121.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@133121.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@133121.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@133135.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@133135.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@133135.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@133135.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@133135.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@133135.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@133149.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@133149.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@133149.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@133149.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@133149.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@133149.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@133163.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@133163.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@133163.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@133163.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@133163.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@133163.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@133177.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@133177.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@133177.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@133177.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@133177.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@133177.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@133191.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@133191.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@133191.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@133191.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@133191.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@133191.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@133205.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@133205.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@133205.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@133205.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@133205.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@133205.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@133219.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@133219.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@133219.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@133219.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@133219.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@133219.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@133233.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@133233.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@133233.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@133233.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@133233.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@133233.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@133247.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@133247.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@133247.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@133247.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@133247.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@133247.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@133261.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@133261.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@133261.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@133261.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@133261.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@133261.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@133275.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@133275.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@133275.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@133275.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@133275.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@133275.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@133289.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@133289.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@133289.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@133289.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@133289.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@133289.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@133303.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@133303.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@133303.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@133303.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@133303.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@133303.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@133317.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@133317.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@133317.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@133317.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@133317.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@133317.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@133331.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@133331.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@133331.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@133331.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@133331.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@133331.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@133345.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@133345.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@133345.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@133345.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@133345.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@133345.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@133359.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@133359.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@133359.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@133359.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@133359.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@133359.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@133373.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@133373.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@133373.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@133373.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@133373.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@133373.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@133387.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@133387.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@133387.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@133387.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@133387.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@133387.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@133401.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@133401.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@133401.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@133401.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@133401.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@133401.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@133415.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@133415.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@133415.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@133415.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@133415.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@133415.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@133429.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@133429.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@133429.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@133429.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@133429.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@133429.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@133443.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@133443.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@133443.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@133443.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@133443.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@133443.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@133457.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@133457.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@133457.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@133457.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@133457.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@133457.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@133471.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@133471.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@133471.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@133471.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@133471.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@133471.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@133485.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@133485.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@133485.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@133485.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@133485.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@133485.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@133499.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@133499.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@133499.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@133499.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@133499.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@133499.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@133513.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@133513.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@133513.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@133513.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@133513.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@133513.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@133527.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@133527.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@133527.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@133527.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@133527.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@133527.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@133541.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@133541.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@133541.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@133541.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@133541.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@133541.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@133555.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@133555.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@133555.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@133555.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@133555.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@133555.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@133569.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@133569.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@133569.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@133569.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@133569.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@133569.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@133583.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@133583.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@133583.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@133583.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@133583.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@133583.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@133597.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@133597.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@133597.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@133597.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@133597.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@133597.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@133611.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@133611.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@133611.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@133611.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@133611.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@133611.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@133625.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@133625.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@133625.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@133625.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@133625.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@133625.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@133639.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@133639.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@133639.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@133639.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@133639.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@133639.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@133653.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@133653.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@133653.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@133653.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@133653.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@133653.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@133667.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@133667.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@133667.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@133667.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@133667.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@133667.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@133681.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@133681.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@133681.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@133681.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@133681.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@133681.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@133695.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@133695.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@133709.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@133709.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@133709.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@133709.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@133709.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@133709.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@133723.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@133723.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@133723.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@133723.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@133723.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@133723.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@133737.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@133737.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@133737.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@133737.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@133737.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@133737.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@133751.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@133751.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@133751.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@133751.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@133751.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@133751.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@133765.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@133765.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@133765.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@133765.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@133765.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@133765.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@133779.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@133779.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@133779.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@133779.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@133779.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@133779.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@133793.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@133793.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@133793.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@133793.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@133793.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@133793.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@133807.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@133807.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@133807.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@133807.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@133807.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@133807.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@133821.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@133821.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@133821.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@133821.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@133821.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@133821.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@133835.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@133835.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@133835.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@133835.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@133835.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@133835.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@133849.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@133849.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@133849.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@133849.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@133849.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@133849.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@133863.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@133863.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@133863.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@133863.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@133863.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@133863.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@133877.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@133877.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@133877.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@133877.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@133877.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@133877.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@133891.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@133891.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@133891.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@133891.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@133891.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@133891.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@133905.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@133905.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@133905.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@133905.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@133905.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@133905.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@133919.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@133919.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@133919.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@133919.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@133919.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@133919.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@133933.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@133933.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@133933.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@133933.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@133933.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@133933.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@133947.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@133947.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@133947.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@133947.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@133947.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@133947.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@133961.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@133961.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@133961.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@133961.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@133961.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@133961.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@133975.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@133975.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@133975.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@133975.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@133975.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@133975.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@133989.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@133989.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@133989.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@133989.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@133989.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@133989.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@134003.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@134003.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@134003.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@134003.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@134003.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@134003.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@134017.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@134017.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@134017.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@134017.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@134017.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@134017.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@134031.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@134031.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@134031.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@134031.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@134031.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@134031.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@134045.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@134045.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@134045.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@134045.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@134045.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@134045.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@134059.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@134059.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@134059.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@134059.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@134059.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@134059.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@134073.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@134073.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@134073.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@134073.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@134073.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@134073.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@134087.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@134087.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@134087.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@134087.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@134087.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@134087.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@134101.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@134101.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@134101.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@134101.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@134101.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@134101.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@134115.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@134115.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@134115.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@134115.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@134115.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@134115.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@134129.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@134129.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@134129.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@134129.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@134129.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@134129.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@134143.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@134143.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@134143.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@134143.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@134143.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@134143.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@134157.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@134157.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@134157.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@134157.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@134157.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@134157.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@134171.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@134171.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@134171.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@134171.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@134171.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@134171.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@134185.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@134185.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@134185.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@134185.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@134185.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@134185.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@134199.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@134199.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@134199.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@134199.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@134199.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@134199.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@134213.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@134213.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@134213.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@134213.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@134213.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@134213.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@134227.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@134227.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@134227.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@134227.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@134227.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@134227.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@134241.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@134241.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@134241.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@134241.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@134241.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@134241.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@134255.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@134255.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@134255.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@134255.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@134255.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@134255.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@134269.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@134269.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@134269.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@134269.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@134269.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@134269.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@134283.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@134283.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@134283.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@134283.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@134283.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@134283.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@134297.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@134297.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@134297.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@134297.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@134297.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@134297.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@134311.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@134311.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@134311.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@134311.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@134311.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@134311.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@134325.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@134325.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@134325.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@134325.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@134325.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@134325.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@134339.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@134339.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@134339.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@134339.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@134339.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@134339.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@134353.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@134353.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@134353.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@134353.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@134353.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@134353.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@134367.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@134367.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@134367.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@134367.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@134367.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@134367.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@134381.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@134381.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@134381.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@134381.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@134381.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@134381.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@134395.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@134395.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@134395.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@134395.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@134395.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@134395.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@134409.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@134409.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@134409.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@134409.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@134409.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@134409.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@134423.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@134423.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@134423.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@134423.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@134423.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@134423.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@134437.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@134437.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@134437.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@134437.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@134437.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@134437.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@134451.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@134451.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@134451.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@134451.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@134451.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@134451.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@134465.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@134465.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@134465.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@134465.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@134465.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@134465.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@134479.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@134479.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@134479.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@134479.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@134479.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@134479.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@134493.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@134493.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@134493.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@134493.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@134493.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@134493.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@134507.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@134507.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@134507.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@134507.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@134507.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@134507.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@134521.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@134521.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@134521.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@134521.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@134521.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@134521.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@134535.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@134535.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@134535.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@134535.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@134535.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@134535.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@134549.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@134549.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@134549.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@134549.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@134549.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@134549.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@134563.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@134563.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@134563.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@134563.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@134563.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@134563.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@134577.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@134577.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@134577.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@134577.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@134577.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@134577.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@134591.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@134591.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@134591.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@134591.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@134591.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@134591.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@134605.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@134605.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@134605.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@134605.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@134605.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@134605.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@134619.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@134619.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@134619.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@134619.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@134619.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@134619.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@134633.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@134633.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@134633.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@134633.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@134633.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@134633.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@134647.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@134647.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@134647.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@134647.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@134647.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@134647.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@134661.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@134661.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@134661.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@134661.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@134661.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@134661.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@134675.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@134675.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@134675.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@134675.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@134675.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@134675.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@134689.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@134689.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@134689.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@134689.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@134689.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@134689.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@134703.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@134703.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@134703.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@134703.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@134703.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@134703.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@134717.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@134717.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@134717.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@134717.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@134717.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@134717.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@134731.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@134731.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@134731.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@134731.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@134731.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@134731.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@134745.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@134745.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@134745.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@134745.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@134745.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@134745.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@134759.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@134759.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@134759.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@134759.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@134759.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@134759.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@134773.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@134773.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@134773.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@134773.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@134773.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@134773.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@134787.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@134787.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@134787.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@134787.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@134787.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@134787.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@134801.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@134801.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@134801.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@134801.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@134801.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@134801.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@134815.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@134815.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@134815.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@134815.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@134815.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@134815.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@134829.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@134829.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@134829.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@134829.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@134829.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@134829.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@134843.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@134843.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@134843.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@134843.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@134843.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@134843.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@134857.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@134857.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@134857.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@134857.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@134857.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@134857.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@134871.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@134871.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@134871.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@134871.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@134871.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@134871.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@134885.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@134885.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@134885.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@134885.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@134885.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@134885.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@134899.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@134899.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@134899.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@134899.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@134899.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@134899.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@134913.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@134913.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@134913.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@127875.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@127887.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@127888.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@127906.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@127918.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@127930.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@127931.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@127872.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@127884.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@127903.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@127915.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@127927.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@127941.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@127955.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@127969.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@127983.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@127997.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@128011.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@128025.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@128039.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@128053.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@128067.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@128081.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@128095.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@128109.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@128123.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@128137.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@128151.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@128165.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@128179.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@128193.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@128207.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@128221.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@128235.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@128249.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@128263.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@128277.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@128291.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@128305.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@128319.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@128333.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@128347.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@128361.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@128375.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@128389.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@128403.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@128417.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@128431.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@128445.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@128459.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@128473.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@128487.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@128501.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@128515.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@128529.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@128543.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@128557.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@128571.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@128585.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@128599.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@128613.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@128627.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@128641.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@128655.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@128669.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@128683.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@128697.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@128711.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@128725.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@128739.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@128753.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@128767.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@128781.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@128795.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@128809.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@128823.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@128837.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@128851.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@128865.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@128879.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@128893.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@128907.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@128921.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@128935.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@128949.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@128963.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@128977.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@128991.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@129005.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@129019.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@129033.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@129047.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@129061.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@129075.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@129089.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@129103.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@129117.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@129131.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@129145.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@129159.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@129173.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@129187.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@129201.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@129215.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@129229.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@129243.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@129257.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@129271.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@129285.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@129299.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@129313.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@129327.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@129341.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@129355.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@129369.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@129383.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@129397.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@129411.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@129425.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@129439.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@129453.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@129467.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@129481.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@129495.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@129509.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@129523.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@129537.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@129551.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@129565.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@129579.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@129593.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@129607.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@129621.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@129635.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@129649.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@129663.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@129677.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@129691.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@129705.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@129719.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@129733.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@129747.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@129761.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@129775.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@129789.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@129803.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@129817.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@129831.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@129845.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@129859.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@129873.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@129887.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@129901.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@129915.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@129929.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@129943.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@129957.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@129971.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@129985.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@129999.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@130013.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@130027.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@130041.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@130055.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@130069.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@130083.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@130097.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@130111.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@130125.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@130139.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@130153.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@130167.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@130181.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@130195.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@130209.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@130223.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@130237.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@130251.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@130265.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@130279.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@130293.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@130307.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@130321.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@130335.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@130349.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@130363.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@130377.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@130391.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@130405.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@130419.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@130433.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@130447.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@130461.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@130475.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@130489.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@130503.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@130517.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@130531.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@130545.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@130559.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@130573.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@130587.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@130601.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@130615.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@130629.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@130643.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@130657.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@130671.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@130685.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@130699.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@130713.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@130727.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@130741.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@130755.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@130769.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@130783.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@130797.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@130811.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@130825.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@130839.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@130853.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@130867.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@130881.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@130895.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@130909.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@130923.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@130937.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@130951.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@130965.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@130979.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@130993.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@131007.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@131021.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@131035.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@131049.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@131063.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@131077.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@131091.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@131105.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@131119.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@131133.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@131147.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@131161.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@131175.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@131189.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@131203.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@131217.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@131231.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@131245.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@131259.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@131273.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@131287.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@131301.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@131315.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@131329.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@131343.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@131357.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@131371.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@131385.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@131399.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@131413.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@131427.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@131441.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@131455.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@131469.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@131483.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@131497.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@131511.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@131525.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@131539.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@131553.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@131567.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@131581.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@131595.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@131609.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@131623.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@131637.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@131651.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@131665.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@131679.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@131693.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@131707.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@131721.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@131735.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@131749.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@131763.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@131777.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@131791.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@131805.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@131819.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@131833.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@131847.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@131861.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@131875.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@131889.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@131903.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@131917.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@131931.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@131945.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@131959.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@131973.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@131987.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@132001.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@132015.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@132029.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@132043.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@132057.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@132071.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@132085.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@132099.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@132113.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@132127.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@132141.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@132155.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@132169.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@132183.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@132197.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@132211.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@132225.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@132239.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@132253.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@132267.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@132281.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@132295.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@132309.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@132323.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@132337.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@132351.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@132365.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@132379.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@132393.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@132407.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@132421.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@132435.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@132449.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@132463.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@132477.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@132491.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@132505.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@132519.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@132533.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@132547.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@132561.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@132575.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@132589.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@132603.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@132617.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@132631.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@132645.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@132659.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@132673.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@132687.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@132701.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@132715.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@132729.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@132743.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@132757.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@132771.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@132785.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@132799.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@132813.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@132827.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@132841.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@132855.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@132869.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@132883.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@132897.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@132911.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@132925.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@132939.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@132953.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@132967.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@132981.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@132995.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@133009.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@133023.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@133037.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@133051.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@133065.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@133079.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@133093.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@133107.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@133121.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@133135.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@133149.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@133163.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@133177.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@133191.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@133205.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@133219.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@133233.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@133247.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@133261.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@133275.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@133289.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@133303.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@133317.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@133331.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@133345.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@133359.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@133373.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@133387.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@133401.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@133415.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@133429.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@133443.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@133457.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@133471.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@133485.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@133499.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@133513.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@133527.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@133541.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@133555.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@133569.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@133583.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@133597.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@133611.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@133625.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@133639.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@133653.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@133667.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@133681.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@133695.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@133709.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@133723.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@133737.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@133751.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@133765.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@133779.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@133793.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@133807.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@133821.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@133835.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@133849.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@133863.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@133877.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@133891.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@133905.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@133919.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@133933.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@133947.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@133961.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@133975.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@133989.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@134003.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@134017.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@134031.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@134045.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@134059.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@134073.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@134087.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@134101.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@134115.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@134129.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@134143.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@134157.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@134171.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@134185.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@134199.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@134213.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@134227.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@134241.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@134255.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@134269.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@134283.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@134297.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@134311.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@134325.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@134339.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@134353.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@134367.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@134381.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@134395.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@134409.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@134423.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@134437.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@134451.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@134465.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@134479.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@134493.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@134507.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@134521.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@134535.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@134549.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@134563.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@134577.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@134591.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@134605.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@134619.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@134633.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@134647.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@134661.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@134675.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@134689.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@134703.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@134717.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@134731.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@134745.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@134759.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@134773.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@134787.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@134801.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@134815.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@134829.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@134843.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@134857.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@134871.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@134885.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@134899.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@134913.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@127875.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@127887.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@127888.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@127906.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@127918.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@127930.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@127931.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@135924.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@135930.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@135931.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@135932.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@135933.4]
  assign regs_0_clock = clock; // @[:@127873.4]
  assign regs_0_reset = reset; // @[:@127874.4 RegFile.scala 82:16:@127880.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@127878.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@127882.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@127877.4]
  assign regs_1_clock = clock; // @[:@127885.4]
  assign regs_1_reset = reset; // @[:@127886.4 RegFile.scala 70:16:@127898.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@127896.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@127901.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@127892.4]
  assign regs_2_clock = clock; // @[:@127904.4]
  assign regs_2_reset = reset; // @[:@127905.4 RegFile.scala 82:16:@127911.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@127909.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@127913.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@127908.4]
  assign regs_3_clock = clock; // @[:@127916.4]
  assign regs_3_reset = reset; // @[:@127917.4 RegFile.scala 82:16:@127923.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@127921.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@127925.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@127920.4]
  assign regs_4_clock = clock; // @[:@127928.4]
  assign regs_4_reset = io_reset; // @[:@127929.4 RegFile.scala 76:16:@127936.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@127935.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@127939.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@127933.4]
  assign regs_5_clock = clock; // @[:@127942.4]
  assign regs_5_reset = io_reset; // @[:@127943.4 RegFile.scala 76:16:@127950.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@127949.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@127953.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@127947.4]
  assign regs_6_clock = clock; // @[:@127956.4]
  assign regs_6_reset = io_reset; // @[:@127957.4 RegFile.scala 76:16:@127964.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@127963.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@127967.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@127961.4]
  assign regs_7_clock = clock; // @[:@127970.4]
  assign regs_7_reset = io_reset; // @[:@127971.4 RegFile.scala 76:16:@127978.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@127977.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@127981.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@127975.4]
  assign regs_8_clock = clock; // @[:@127984.4]
  assign regs_8_reset = io_reset; // @[:@127985.4 RegFile.scala 76:16:@127992.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@127991.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@127995.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@127989.4]
  assign regs_9_clock = clock; // @[:@127998.4]
  assign regs_9_reset = io_reset; // @[:@127999.4 RegFile.scala 76:16:@128006.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@128005.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@128009.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@128003.4]
  assign regs_10_clock = clock; // @[:@128012.4]
  assign regs_10_reset = io_reset; // @[:@128013.4 RegFile.scala 76:16:@128020.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@128019.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@128023.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@128017.4]
  assign regs_11_clock = clock; // @[:@128026.4]
  assign regs_11_reset = io_reset; // @[:@128027.4 RegFile.scala 76:16:@128034.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@128033.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@128037.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@128031.4]
  assign regs_12_clock = clock; // @[:@128040.4]
  assign regs_12_reset = io_reset; // @[:@128041.4 RegFile.scala 76:16:@128048.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@128047.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@128051.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@128045.4]
  assign regs_13_clock = clock; // @[:@128054.4]
  assign regs_13_reset = io_reset; // @[:@128055.4 RegFile.scala 76:16:@128062.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@128061.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@128065.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@128059.4]
  assign regs_14_clock = clock; // @[:@128068.4]
  assign regs_14_reset = io_reset; // @[:@128069.4 RegFile.scala 76:16:@128076.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@128075.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@128079.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@128073.4]
  assign regs_15_clock = clock; // @[:@128082.4]
  assign regs_15_reset = io_reset; // @[:@128083.4 RegFile.scala 76:16:@128090.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@128089.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@128093.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@128087.4]
  assign regs_16_clock = clock; // @[:@128096.4]
  assign regs_16_reset = io_reset; // @[:@128097.4 RegFile.scala 76:16:@128104.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@128103.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@128107.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@128101.4]
  assign regs_17_clock = clock; // @[:@128110.4]
  assign regs_17_reset = io_reset; // @[:@128111.4 RegFile.scala 76:16:@128118.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@128117.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@128121.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@128115.4]
  assign regs_18_clock = clock; // @[:@128124.4]
  assign regs_18_reset = io_reset; // @[:@128125.4 RegFile.scala 76:16:@128132.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@128131.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@128135.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@128129.4]
  assign regs_19_clock = clock; // @[:@128138.4]
  assign regs_19_reset = io_reset; // @[:@128139.4 RegFile.scala 76:16:@128146.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@128145.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@128149.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@128143.4]
  assign regs_20_clock = clock; // @[:@128152.4]
  assign regs_20_reset = io_reset; // @[:@128153.4 RegFile.scala 76:16:@128160.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@128159.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@128163.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@128157.4]
  assign regs_21_clock = clock; // @[:@128166.4]
  assign regs_21_reset = io_reset; // @[:@128167.4 RegFile.scala 76:16:@128174.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@128173.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@128177.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@128171.4]
  assign regs_22_clock = clock; // @[:@128180.4]
  assign regs_22_reset = io_reset; // @[:@128181.4 RegFile.scala 76:16:@128188.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@128187.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@128191.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@128185.4]
  assign regs_23_clock = clock; // @[:@128194.4]
  assign regs_23_reset = io_reset; // @[:@128195.4 RegFile.scala 76:16:@128202.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@128201.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@128205.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@128199.4]
  assign regs_24_clock = clock; // @[:@128208.4]
  assign regs_24_reset = io_reset; // @[:@128209.4 RegFile.scala 76:16:@128216.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@128215.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@128219.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@128213.4]
  assign regs_25_clock = clock; // @[:@128222.4]
  assign regs_25_reset = io_reset; // @[:@128223.4 RegFile.scala 76:16:@128230.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@128229.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@128233.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@128227.4]
  assign regs_26_clock = clock; // @[:@128236.4]
  assign regs_26_reset = io_reset; // @[:@128237.4 RegFile.scala 76:16:@128244.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@128243.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@128247.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@128241.4]
  assign regs_27_clock = clock; // @[:@128250.4]
  assign regs_27_reset = io_reset; // @[:@128251.4 RegFile.scala 76:16:@128258.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@128257.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@128261.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@128255.4]
  assign regs_28_clock = clock; // @[:@128264.4]
  assign regs_28_reset = io_reset; // @[:@128265.4 RegFile.scala 76:16:@128272.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@128271.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@128275.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@128269.4]
  assign regs_29_clock = clock; // @[:@128278.4]
  assign regs_29_reset = io_reset; // @[:@128279.4 RegFile.scala 76:16:@128286.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@128285.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@128289.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@128283.4]
  assign regs_30_clock = clock; // @[:@128292.4]
  assign regs_30_reset = io_reset; // @[:@128293.4 RegFile.scala 76:16:@128300.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@128299.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@128303.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@128297.4]
  assign regs_31_clock = clock; // @[:@128306.4]
  assign regs_31_reset = io_reset; // @[:@128307.4 RegFile.scala 76:16:@128314.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@128313.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@128317.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@128311.4]
  assign regs_32_clock = clock; // @[:@128320.4]
  assign regs_32_reset = io_reset; // @[:@128321.4 RegFile.scala 76:16:@128328.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@128327.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@128331.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@128325.4]
  assign regs_33_clock = clock; // @[:@128334.4]
  assign regs_33_reset = io_reset; // @[:@128335.4 RegFile.scala 76:16:@128342.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@128341.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@128345.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@128339.4]
  assign regs_34_clock = clock; // @[:@128348.4]
  assign regs_34_reset = io_reset; // @[:@128349.4 RegFile.scala 76:16:@128356.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@128355.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@128359.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@128353.4]
  assign regs_35_clock = clock; // @[:@128362.4]
  assign regs_35_reset = io_reset; // @[:@128363.4 RegFile.scala 76:16:@128370.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@128369.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@128373.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@128367.4]
  assign regs_36_clock = clock; // @[:@128376.4]
  assign regs_36_reset = io_reset; // @[:@128377.4 RegFile.scala 76:16:@128384.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@128383.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@128387.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@128381.4]
  assign regs_37_clock = clock; // @[:@128390.4]
  assign regs_37_reset = io_reset; // @[:@128391.4 RegFile.scala 76:16:@128398.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@128397.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@128401.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@128395.4]
  assign regs_38_clock = clock; // @[:@128404.4]
  assign regs_38_reset = io_reset; // @[:@128405.4 RegFile.scala 76:16:@128412.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@128411.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@128415.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@128409.4]
  assign regs_39_clock = clock; // @[:@128418.4]
  assign regs_39_reset = io_reset; // @[:@128419.4 RegFile.scala 76:16:@128426.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@128425.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@128429.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@128423.4]
  assign regs_40_clock = clock; // @[:@128432.4]
  assign regs_40_reset = io_reset; // @[:@128433.4 RegFile.scala 76:16:@128440.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@128439.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@128443.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@128437.4]
  assign regs_41_clock = clock; // @[:@128446.4]
  assign regs_41_reset = io_reset; // @[:@128447.4 RegFile.scala 76:16:@128454.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@128453.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@128457.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@128451.4]
  assign regs_42_clock = clock; // @[:@128460.4]
  assign regs_42_reset = io_reset; // @[:@128461.4 RegFile.scala 76:16:@128468.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@128467.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@128471.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@128465.4]
  assign regs_43_clock = clock; // @[:@128474.4]
  assign regs_43_reset = io_reset; // @[:@128475.4 RegFile.scala 76:16:@128482.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@128481.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@128485.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@128479.4]
  assign regs_44_clock = clock; // @[:@128488.4]
  assign regs_44_reset = io_reset; // @[:@128489.4 RegFile.scala 76:16:@128496.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@128495.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@128499.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@128493.4]
  assign regs_45_clock = clock; // @[:@128502.4]
  assign regs_45_reset = io_reset; // @[:@128503.4 RegFile.scala 76:16:@128510.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@128509.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@128513.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@128507.4]
  assign regs_46_clock = clock; // @[:@128516.4]
  assign regs_46_reset = io_reset; // @[:@128517.4 RegFile.scala 76:16:@128524.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@128523.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@128527.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@128521.4]
  assign regs_47_clock = clock; // @[:@128530.4]
  assign regs_47_reset = io_reset; // @[:@128531.4 RegFile.scala 76:16:@128538.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@128537.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@128541.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@128535.4]
  assign regs_48_clock = clock; // @[:@128544.4]
  assign regs_48_reset = io_reset; // @[:@128545.4 RegFile.scala 76:16:@128552.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@128551.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@128555.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@128549.4]
  assign regs_49_clock = clock; // @[:@128558.4]
  assign regs_49_reset = io_reset; // @[:@128559.4 RegFile.scala 76:16:@128566.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@128565.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@128569.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@128563.4]
  assign regs_50_clock = clock; // @[:@128572.4]
  assign regs_50_reset = io_reset; // @[:@128573.4 RegFile.scala 76:16:@128580.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@128579.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@128583.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@128577.4]
  assign regs_51_clock = clock; // @[:@128586.4]
  assign regs_51_reset = io_reset; // @[:@128587.4 RegFile.scala 76:16:@128594.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@128593.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@128597.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@128591.4]
  assign regs_52_clock = clock; // @[:@128600.4]
  assign regs_52_reset = io_reset; // @[:@128601.4 RegFile.scala 76:16:@128608.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@128607.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@128611.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@128605.4]
  assign regs_53_clock = clock; // @[:@128614.4]
  assign regs_53_reset = io_reset; // @[:@128615.4 RegFile.scala 76:16:@128622.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@128621.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@128625.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@128619.4]
  assign regs_54_clock = clock; // @[:@128628.4]
  assign regs_54_reset = io_reset; // @[:@128629.4 RegFile.scala 76:16:@128636.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@128635.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@128639.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@128633.4]
  assign regs_55_clock = clock; // @[:@128642.4]
  assign regs_55_reset = io_reset; // @[:@128643.4 RegFile.scala 76:16:@128650.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@128649.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@128653.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@128647.4]
  assign regs_56_clock = clock; // @[:@128656.4]
  assign regs_56_reset = io_reset; // @[:@128657.4 RegFile.scala 76:16:@128664.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@128663.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@128667.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@128661.4]
  assign regs_57_clock = clock; // @[:@128670.4]
  assign regs_57_reset = io_reset; // @[:@128671.4 RegFile.scala 76:16:@128678.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@128677.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@128681.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@128675.4]
  assign regs_58_clock = clock; // @[:@128684.4]
  assign regs_58_reset = io_reset; // @[:@128685.4 RegFile.scala 76:16:@128692.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@128691.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@128695.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@128689.4]
  assign regs_59_clock = clock; // @[:@128698.4]
  assign regs_59_reset = io_reset; // @[:@128699.4 RegFile.scala 76:16:@128706.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@128705.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@128709.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@128703.4]
  assign regs_60_clock = clock; // @[:@128712.4]
  assign regs_60_reset = io_reset; // @[:@128713.4 RegFile.scala 76:16:@128720.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@128719.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@128723.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@128717.4]
  assign regs_61_clock = clock; // @[:@128726.4]
  assign regs_61_reset = io_reset; // @[:@128727.4 RegFile.scala 76:16:@128734.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@128733.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@128737.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@128731.4]
  assign regs_62_clock = clock; // @[:@128740.4]
  assign regs_62_reset = io_reset; // @[:@128741.4 RegFile.scala 76:16:@128748.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@128747.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@128751.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@128745.4]
  assign regs_63_clock = clock; // @[:@128754.4]
  assign regs_63_reset = io_reset; // @[:@128755.4 RegFile.scala 76:16:@128762.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@128761.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@128765.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@128759.4]
  assign regs_64_clock = clock; // @[:@128768.4]
  assign regs_64_reset = io_reset; // @[:@128769.4 RegFile.scala 76:16:@128776.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@128775.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@128779.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@128773.4]
  assign regs_65_clock = clock; // @[:@128782.4]
  assign regs_65_reset = io_reset; // @[:@128783.4 RegFile.scala 76:16:@128790.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@128789.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@128793.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@128787.4]
  assign regs_66_clock = clock; // @[:@128796.4]
  assign regs_66_reset = io_reset; // @[:@128797.4 RegFile.scala 76:16:@128804.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@128803.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@128807.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@128801.4]
  assign regs_67_clock = clock; // @[:@128810.4]
  assign regs_67_reset = io_reset; // @[:@128811.4 RegFile.scala 76:16:@128818.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@128817.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@128821.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@128815.4]
  assign regs_68_clock = clock; // @[:@128824.4]
  assign regs_68_reset = io_reset; // @[:@128825.4 RegFile.scala 76:16:@128832.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@128831.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@128835.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@128829.4]
  assign regs_69_clock = clock; // @[:@128838.4]
  assign regs_69_reset = io_reset; // @[:@128839.4 RegFile.scala 76:16:@128846.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@128845.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@128849.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@128843.4]
  assign regs_70_clock = clock; // @[:@128852.4]
  assign regs_70_reset = io_reset; // @[:@128853.4 RegFile.scala 76:16:@128860.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@128859.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@128863.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@128857.4]
  assign regs_71_clock = clock; // @[:@128866.4]
  assign regs_71_reset = io_reset; // @[:@128867.4 RegFile.scala 76:16:@128874.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@128873.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@128877.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@128871.4]
  assign regs_72_clock = clock; // @[:@128880.4]
  assign regs_72_reset = io_reset; // @[:@128881.4 RegFile.scala 76:16:@128888.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@128887.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@128891.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@128885.4]
  assign regs_73_clock = clock; // @[:@128894.4]
  assign regs_73_reset = io_reset; // @[:@128895.4 RegFile.scala 76:16:@128902.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@128901.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@128905.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@128899.4]
  assign regs_74_clock = clock; // @[:@128908.4]
  assign regs_74_reset = io_reset; // @[:@128909.4 RegFile.scala 76:16:@128916.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@128915.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@128919.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@128913.4]
  assign regs_75_clock = clock; // @[:@128922.4]
  assign regs_75_reset = io_reset; // @[:@128923.4 RegFile.scala 76:16:@128930.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@128929.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@128933.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@128927.4]
  assign regs_76_clock = clock; // @[:@128936.4]
  assign regs_76_reset = io_reset; // @[:@128937.4 RegFile.scala 76:16:@128944.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@128943.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@128947.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@128941.4]
  assign regs_77_clock = clock; // @[:@128950.4]
  assign regs_77_reset = io_reset; // @[:@128951.4 RegFile.scala 76:16:@128958.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@128957.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@128961.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@128955.4]
  assign regs_78_clock = clock; // @[:@128964.4]
  assign regs_78_reset = io_reset; // @[:@128965.4 RegFile.scala 76:16:@128972.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@128971.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@128975.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@128969.4]
  assign regs_79_clock = clock; // @[:@128978.4]
  assign regs_79_reset = io_reset; // @[:@128979.4 RegFile.scala 76:16:@128986.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@128985.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@128989.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@128983.4]
  assign regs_80_clock = clock; // @[:@128992.4]
  assign regs_80_reset = io_reset; // @[:@128993.4 RegFile.scala 76:16:@129000.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@128999.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@129003.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@128997.4]
  assign regs_81_clock = clock; // @[:@129006.4]
  assign regs_81_reset = io_reset; // @[:@129007.4 RegFile.scala 76:16:@129014.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@129013.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@129017.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@129011.4]
  assign regs_82_clock = clock; // @[:@129020.4]
  assign regs_82_reset = io_reset; // @[:@129021.4 RegFile.scala 76:16:@129028.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@129027.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@129031.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@129025.4]
  assign regs_83_clock = clock; // @[:@129034.4]
  assign regs_83_reset = io_reset; // @[:@129035.4 RegFile.scala 76:16:@129042.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@129041.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@129045.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@129039.4]
  assign regs_84_clock = clock; // @[:@129048.4]
  assign regs_84_reset = io_reset; // @[:@129049.4 RegFile.scala 76:16:@129056.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@129055.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@129059.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@129053.4]
  assign regs_85_clock = clock; // @[:@129062.4]
  assign regs_85_reset = io_reset; // @[:@129063.4 RegFile.scala 76:16:@129070.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@129069.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@129073.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@129067.4]
  assign regs_86_clock = clock; // @[:@129076.4]
  assign regs_86_reset = io_reset; // @[:@129077.4 RegFile.scala 76:16:@129084.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@129083.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@129087.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@129081.4]
  assign regs_87_clock = clock; // @[:@129090.4]
  assign regs_87_reset = io_reset; // @[:@129091.4 RegFile.scala 76:16:@129098.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@129097.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@129101.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@129095.4]
  assign regs_88_clock = clock; // @[:@129104.4]
  assign regs_88_reset = io_reset; // @[:@129105.4 RegFile.scala 76:16:@129112.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@129111.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@129115.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@129109.4]
  assign regs_89_clock = clock; // @[:@129118.4]
  assign regs_89_reset = io_reset; // @[:@129119.4 RegFile.scala 76:16:@129126.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@129125.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@129129.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@129123.4]
  assign regs_90_clock = clock; // @[:@129132.4]
  assign regs_90_reset = io_reset; // @[:@129133.4 RegFile.scala 76:16:@129140.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@129139.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@129143.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@129137.4]
  assign regs_91_clock = clock; // @[:@129146.4]
  assign regs_91_reset = io_reset; // @[:@129147.4 RegFile.scala 76:16:@129154.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@129153.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@129157.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@129151.4]
  assign regs_92_clock = clock; // @[:@129160.4]
  assign regs_92_reset = io_reset; // @[:@129161.4 RegFile.scala 76:16:@129168.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@129167.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@129171.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@129165.4]
  assign regs_93_clock = clock; // @[:@129174.4]
  assign regs_93_reset = io_reset; // @[:@129175.4 RegFile.scala 76:16:@129182.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@129181.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@129185.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@129179.4]
  assign regs_94_clock = clock; // @[:@129188.4]
  assign regs_94_reset = io_reset; // @[:@129189.4 RegFile.scala 76:16:@129196.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@129195.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@129199.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@129193.4]
  assign regs_95_clock = clock; // @[:@129202.4]
  assign regs_95_reset = io_reset; // @[:@129203.4 RegFile.scala 76:16:@129210.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@129209.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@129213.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@129207.4]
  assign regs_96_clock = clock; // @[:@129216.4]
  assign regs_96_reset = io_reset; // @[:@129217.4 RegFile.scala 76:16:@129224.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@129223.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@129227.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@129221.4]
  assign regs_97_clock = clock; // @[:@129230.4]
  assign regs_97_reset = io_reset; // @[:@129231.4 RegFile.scala 76:16:@129238.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@129237.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@129241.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@129235.4]
  assign regs_98_clock = clock; // @[:@129244.4]
  assign regs_98_reset = io_reset; // @[:@129245.4 RegFile.scala 76:16:@129252.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@129251.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@129255.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@129249.4]
  assign regs_99_clock = clock; // @[:@129258.4]
  assign regs_99_reset = io_reset; // @[:@129259.4 RegFile.scala 76:16:@129266.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@129265.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@129269.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@129263.4]
  assign regs_100_clock = clock; // @[:@129272.4]
  assign regs_100_reset = io_reset; // @[:@129273.4 RegFile.scala 76:16:@129280.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@129279.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@129283.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@129277.4]
  assign regs_101_clock = clock; // @[:@129286.4]
  assign regs_101_reset = io_reset; // @[:@129287.4 RegFile.scala 76:16:@129294.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@129293.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@129297.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@129291.4]
  assign regs_102_clock = clock; // @[:@129300.4]
  assign regs_102_reset = io_reset; // @[:@129301.4 RegFile.scala 76:16:@129308.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@129307.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@129311.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@129305.4]
  assign regs_103_clock = clock; // @[:@129314.4]
  assign regs_103_reset = io_reset; // @[:@129315.4 RegFile.scala 76:16:@129322.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@129321.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@129325.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@129319.4]
  assign regs_104_clock = clock; // @[:@129328.4]
  assign regs_104_reset = io_reset; // @[:@129329.4 RegFile.scala 76:16:@129336.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@129335.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@129339.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@129333.4]
  assign regs_105_clock = clock; // @[:@129342.4]
  assign regs_105_reset = io_reset; // @[:@129343.4 RegFile.scala 76:16:@129350.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@129349.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@129353.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@129347.4]
  assign regs_106_clock = clock; // @[:@129356.4]
  assign regs_106_reset = io_reset; // @[:@129357.4 RegFile.scala 76:16:@129364.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@129363.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@129367.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@129361.4]
  assign regs_107_clock = clock; // @[:@129370.4]
  assign regs_107_reset = io_reset; // @[:@129371.4 RegFile.scala 76:16:@129378.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@129377.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@129381.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@129375.4]
  assign regs_108_clock = clock; // @[:@129384.4]
  assign regs_108_reset = io_reset; // @[:@129385.4 RegFile.scala 76:16:@129392.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@129391.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@129395.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@129389.4]
  assign regs_109_clock = clock; // @[:@129398.4]
  assign regs_109_reset = io_reset; // @[:@129399.4 RegFile.scala 76:16:@129406.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@129405.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@129409.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@129403.4]
  assign regs_110_clock = clock; // @[:@129412.4]
  assign regs_110_reset = io_reset; // @[:@129413.4 RegFile.scala 76:16:@129420.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@129419.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@129423.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@129417.4]
  assign regs_111_clock = clock; // @[:@129426.4]
  assign regs_111_reset = io_reset; // @[:@129427.4 RegFile.scala 76:16:@129434.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@129433.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@129437.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@129431.4]
  assign regs_112_clock = clock; // @[:@129440.4]
  assign regs_112_reset = io_reset; // @[:@129441.4 RegFile.scala 76:16:@129448.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@129447.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@129451.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@129445.4]
  assign regs_113_clock = clock; // @[:@129454.4]
  assign regs_113_reset = io_reset; // @[:@129455.4 RegFile.scala 76:16:@129462.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@129461.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@129465.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@129459.4]
  assign regs_114_clock = clock; // @[:@129468.4]
  assign regs_114_reset = io_reset; // @[:@129469.4 RegFile.scala 76:16:@129476.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@129475.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@129479.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@129473.4]
  assign regs_115_clock = clock; // @[:@129482.4]
  assign regs_115_reset = io_reset; // @[:@129483.4 RegFile.scala 76:16:@129490.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@129489.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@129493.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@129487.4]
  assign regs_116_clock = clock; // @[:@129496.4]
  assign regs_116_reset = io_reset; // @[:@129497.4 RegFile.scala 76:16:@129504.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@129503.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@129507.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@129501.4]
  assign regs_117_clock = clock; // @[:@129510.4]
  assign regs_117_reset = io_reset; // @[:@129511.4 RegFile.scala 76:16:@129518.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@129517.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@129521.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@129515.4]
  assign regs_118_clock = clock; // @[:@129524.4]
  assign regs_118_reset = io_reset; // @[:@129525.4 RegFile.scala 76:16:@129532.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@129531.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@129535.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@129529.4]
  assign regs_119_clock = clock; // @[:@129538.4]
  assign regs_119_reset = io_reset; // @[:@129539.4 RegFile.scala 76:16:@129546.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@129545.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@129549.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@129543.4]
  assign regs_120_clock = clock; // @[:@129552.4]
  assign regs_120_reset = io_reset; // @[:@129553.4 RegFile.scala 76:16:@129560.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@129559.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@129563.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@129557.4]
  assign regs_121_clock = clock; // @[:@129566.4]
  assign regs_121_reset = io_reset; // @[:@129567.4 RegFile.scala 76:16:@129574.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@129573.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@129577.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@129571.4]
  assign regs_122_clock = clock; // @[:@129580.4]
  assign regs_122_reset = io_reset; // @[:@129581.4 RegFile.scala 76:16:@129588.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@129587.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@129591.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@129585.4]
  assign regs_123_clock = clock; // @[:@129594.4]
  assign regs_123_reset = io_reset; // @[:@129595.4 RegFile.scala 76:16:@129602.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@129601.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@129605.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@129599.4]
  assign regs_124_clock = clock; // @[:@129608.4]
  assign regs_124_reset = io_reset; // @[:@129609.4 RegFile.scala 76:16:@129616.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@129615.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@129619.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@129613.4]
  assign regs_125_clock = clock; // @[:@129622.4]
  assign regs_125_reset = io_reset; // @[:@129623.4 RegFile.scala 76:16:@129630.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@129629.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@129633.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@129627.4]
  assign regs_126_clock = clock; // @[:@129636.4]
  assign regs_126_reset = io_reset; // @[:@129637.4 RegFile.scala 76:16:@129644.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@129643.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@129647.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@129641.4]
  assign regs_127_clock = clock; // @[:@129650.4]
  assign regs_127_reset = io_reset; // @[:@129651.4 RegFile.scala 76:16:@129658.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@129657.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@129661.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@129655.4]
  assign regs_128_clock = clock; // @[:@129664.4]
  assign regs_128_reset = io_reset; // @[:@129665.4 RegFile.scala 76:16:@129672.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@129671.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@129675.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@129669.4]
  assign regs_129_clock = clock; // @[:@129678.4]
  assign regs_129_reset = io_reset; // @[:@129679.4 RegFile.scala 76:16:@129686.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@129685.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@129689.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@129683.4]
  assign regs_130_clock = clock; // @[:@129692.4]
  assign regs_130_reset = io_reset; // @[:@129693.4 RegFile.scala 76:16:@129700.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@129699.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@129703.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@129697.4]
  assign regs_131_clock = clock; // @[:@129706.4]
  assign regs_131_reset = io_reset; // @[:@129707.4 RegFile.scala 76:16:@129714.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@129713.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@129717.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@129711.4]
  assign regs_132_clock = clock; // @[:@129720.4]
  assign regs_132_reset = io_reset; // @[:@129721.4 RegFile.scala 76:16:@129728.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@129727.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@129731.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@129725.4]
  assign regs_133_clock = clock; // @[:@129734.4]
  assign regs_133_reset = io_reset; // @[:@129735.4 RegFile.scala 76:16:@129742.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@129741.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@129745.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@129739.4]
  assign regs_134_clock = clock; // @[:@129748.4]
  assign regs_134_reset = io_reset; // @[:@129749.4 RegFile.scala 76:16:@129756.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@129755.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@129759.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@129753.4]
  assign regs_135_clock = clock; // @[:@129762.4]
  assign regs_135_reset = io_reset; // @[:@129763.4 RegFile.scala 76:16:@129770.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@129769.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@129773.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@129767.4]
  assign regs_136_clock = clock; // @[:@129776.4]
  assign regs_136_reset = io_reset; // @[:@129777.4 RegFile.scala 76:16:@129784.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@129783.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@129787.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@129781.4]
  assign regs_137_clock = clock; // @[:@129790.4]
  assign regs_137_reset = io_reset; // @[:@129791.4 RegFile.scala 76:16:@129798.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@129797.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@129801.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@129795.4]
  assign regs_138_clock = clock; // @[:@129804.4]
  assign regs_138_reset = io_reset; // @[:@129805.4 RegFile.scala 76:16:@129812.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@129811.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@129815.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@129809.4]
  assign regs_139_clock = clock; // @[:@129818.4]
  assign regs_139_reset = io_reset; // @[:@129819.4 RegFile.scala 76:16:@129826.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@129825.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@129829.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@129823.4]
  assign regs_140_clock = clock; // @[:@129832.4]
  assign regs_140_reset = io_reset; // @[:@129833.4 RegFile.scala 76:16:@129840.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@129839.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@129843.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@129837.4]
  assign regs_141_clock = clock; // @[:@129846.4]
  assign regs_141_reset = io_reset; // @[:@129847.4 RegFile.scala 76:16:@129854.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@129853.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@129857.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@129851.4]
  assign regs_142_clock = clock; // @[:@129860.4]
  assign regs_142_reset = io_reset; // @[:@129861.4 RegFile.scala 76:16:@129868.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@129867.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@129871.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@129865.4]
  assign regs_143_clock = clock; // @[:@129874.4]
  assign regs_143_reset = io_reset; // @[:@129875.4 RegFile.scala 76:16:@129882.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@129881.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@129885.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@129879.4]
  assign regs_144_clock = clock; // @[:@129888.4]
  assign regs_144_reset = io_reset; // @[:@129889.4 RegFile.scala 76:16:@129896.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@129895.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@129899.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@129893.4]
  assign regs_145_clock = clock; // @[:@129902.4]
  assign regs_145_reset = io_reset; // @[:@129903.4 RegFile.scala 76:16:@129910.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@129909.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@129913.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@129907.4]
  assign regs_146_clock = clock; // @[:@129916.4]
  assign regs_146_reset = io_reset; // @[:@129917.4 RegFile.scala 76:16:@129924.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@129923.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@129927.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@129921.4]
  assign regs_147_clock = clock; // @[:@129930.4]
  assign regs_147_reset = io_reset; // @[:@129931.4 RegFile.scala 76:16:@129938.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@129937.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@129941.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@129935.4]
  assign regs_148_clock = clock; // @[:@129944.4]
  assign regs_148_reset = io_reset; // @[:@129945.4 RegFile.scala 76:16:@129952.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@129951.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@129955.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@129949.4]
  assign regs_149_clock = clock; // @[:@129958.4]
  assign regs_149_reset = io_reset; // @[:@129959.4 RegFile.scala 76:16:@129966.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@129965.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@129969.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@129963.4]
  assign regs_150_clock = clock; // @[:@129972.4]
  assign regs_150_reset = io_reset; // @[:@129973.4 RegFile.scala 76:16:@129980.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@129979.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@129983.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@129977.4]
  assign regs_151_clock = clock; // @[:@129986.4]
  assign regs_151_reset = io_reset; // @[:@129987.4 RegFile.scala 76:16:@129994.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@129993.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@129997.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@129991.4]
  assign regs_152_clock = clock; // @[:@130000.4]
  assign regs_152_reset = io_reset; // @[:@130001.4 RegFile.scala 76:16:@130008.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@130007.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@130011.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@130005.4]
  assign regs_153_clock = clock; // @[:@130014.4]
  assign regs_153_reset = io_reset; // @[:@130015.4 RegFile.scala 76:16:@130022.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@130021.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@130025.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@130019.4]
  assign regs_154_clock = clock; // @[:@130028.4]
  assign regs_154_reset = io_reset; // @[:@130029.4 RegFile.scala 76:16:@130036.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@130035.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@130039.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@130033.4]
  assign regs_155_clock = clock; // @[:@130042.4]
  assign regs_155_reset = io_reset; // @[:@130043.4 RegFile.scala 76:16:@130050.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@130049.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@130053.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@130047.4]
  assign regs_156_clock = clock; // @[:@130056.4]
  assign regs_156_reset = io_reset; // @[:@130057.4 RegFile.scala 76:16:@130064.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@130063.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@130067.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@130061.4]
  assign regs_157_clock = clock; // @[:@130070.4]
  assign regs_157_reset = io_reset; // @[:@130071.4 RegFile.scala 76:16:@130078.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@130077.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@130081.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@130075.4]
  assign regs_158_clock = clock; // @[:@130084.4]
  assign regs_158_reset = io_reset; // @[:@130085.4 RegFile.scala 76:16:@130092.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@130091.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@130095.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@130089.4]
  assign regs_159_clock = clock; // @[:@130098.4]
  assign regs_159_reset = io_reset; // @[:@130099.4 RegFile.scala 76:16:@130106.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@130105.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@130109.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@130103.4]
  assign regs_160_clock = clock; // @[:@130112.4]
  assign regs_160_reset = io_reset; // @[:@130113.4 RegFile.scala 76:16:@130120.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@130119.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@130123.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@130117.4]
  assign regs_161_clock = clock; // @[:@130126.4]
  assign regs_161_reset = io_reset; // @[:@130127.4 RegFile.scala 76:16:@130134.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@130133.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@130137.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@130131.4]
  assign regs_162_clock = clock; // @[:@130140.4]
  assign regs_162_reset = io_reset; // @[:@130141.4 RegFile.scala 76:16:@130148.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@130147.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@130151.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@130145.4]
  assign regs_163_clock = clock; // @[:@130154.4]
  assign regs_163_reset = io_reset; // @[:@130155.4 RegFile.scala 76:16:@130162.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@130161.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@130165.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@130159.4]
  assign regs_164_clock = clock; // @[:@130168.4]
  assign regs_164_reset = io_reset; // @[:@130169.4 RegFile.scala 76:16:@130176.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@130175.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@130179.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@130173.4]
  assign regs_165_clock = clock; // @[:@130182.4]
  assign regs_165_reset = io_reset; // @[:@130183.4 RegFile.scala 76:16:@130190.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@130189.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@130193.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@130187.4]
  assign regs_166_clock = clock; // @[:@130196.4]
  assign regs_166_reset = io_reset; // @[:@130197.4 RegFile.scala 76:16:@130204.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@130203.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@130207.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@130201.4]
  assign regs_167_clock = clock; // @[:@130210.4]
  assign regs_167_reset = io_reset; // @[:@130211.4 RegFile.scala 76:16:@130218.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@130217.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@130221.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@130215.4]
  assign regs_168_clock = clock; // @[:@130224.4]
  assign regs_168_reset = io_reset; // @[:@130225.4 RegFile.scala 76:16:@130232.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@130231.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@130235.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@130229.4]
  assign regs_169_clock = clock; // @[:@130238.4]
  assign regs_169_reset = io_reset; // @[:@130239.4 RegFile.scala 76:16:@130246.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@130245.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@130249.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@130243.4]
  assign regs_170_clock = clock; // @[:@130252.4]
  assign regs_170_reset = io_reset; // @[:@130253.4 RegFile.scala 76:16:@130260.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@130259.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@130263.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@130257.4]
  assign regs_171_clock = clock; // @[:@130266.4]
  assign regs_171_reset = io_reset; // @[:@130267.4 RegFile.scala 76:16:@130274.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@130273.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@130277.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@130271.4]
  assign regs_172_clock = clock; // @[:@130280.4]
  assign regs_172_reset = io_reset; // @[:@130281.4 RegFile.scala 76:16:@130288.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@130287.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@130291.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@130285.4]
  assign regs_173_clock = clock; // @[:@130294.4]
  assign regs_173_reset = io_reset; // @[:@130295.4 RegFile.scala 76:16:@130302.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@130301.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@130305.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@130299.4]
  assign regs_174_clock = clock; // @[:@130308.4]
  assign regs_174_reset = io_reset; // @[:@130309.4 RegFile.scala 76:16:@130316.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@130315.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@130319.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@130313.4]
  assign regs_175_clock = clock; // @[:@130322.4]
  assign regs_175_reset = io_reset; // @[:@130323.4 RegFile.scala 76:16:@130330.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@130329.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@130333.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@130327.4]
  assign regs_176_clock = clock; // @[:@130336.4]
  assign regs_176_reset = io_reset; // @[:@130337.4 RegFile.scala 76:16:@130344.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@130343.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@130347.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@130341.4]
  assign regs_177_clock = clock; // @[:@130350.4]
  assign regs_177_reset = io_reset; // @[:@130351.4 RegFile.scala 76:16:@130358.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@130357.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@130361.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@130355.4]
  assign regs_178_clock = clock; // @[:@130364.4]
  assign regs_178_reset = io_reset; // @[:@130365.4 RegFile.scala 76:16:@130372.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@130371.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@130375.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@130369.4]
  assign regs_179_clock = clock; // @[:@130378.4]
  assign regs_179_reset = io_reset; // @[:@130379.4 RegFile.scala 76:16:@130386.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@130385.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@130389.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@130383.4]
  assign regs_180_clock = clock; // @[:@130392.4]
  assign regs_180_reset = io_reset; // @[:@130393.4 RegFile.scala 76:16:@130400.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@130399.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@130403.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@130397.4]
  assign regs_181_clock = clock; // @[:@130406.4]
  assign regs_181_reset = io_reset; // @[:@130407.4 RegFile.scala 76:16:@130414.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@130413.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@130417.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@130411.4]
  assign regs_182_clock = clock; // @[:@130420.4]
  assign regs_182_reset = io_reset; // @[:@130421.4 RegFile.scala 76:16:@130428.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@130427.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@130431.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@130425.4]
  assign regs_183_clock = clock; // @[:@130434.4]
  assign regs_183_reset = io_reset; // @[:@130435.4 RegFile.scala 76:16:@130442.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@130441.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@130445.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@130439.4]
  assign regs_184_clock = clock; // @[:@130448.4]
  assign regs_184_reset = io_reset; // @[:@130449.4 RegFile.scala 76:16:@130456.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@130455.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@130459.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@130453.4]
  assign regs_185_clock = clock; // @[:@130462.4]
  assign regs_185_reset = io_reset; // @[:@130463.4 RegFile.scala 76:16:@130470.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@130469.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@130473.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@130467.4]
  assign regs_186_clock = clock; // @[:@130476.4]
  assign regs_186_reset = io_reset; // @[:@130477.4 RegFile.scala 76:16:@130484.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@130483.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@130487.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@130481.4]
  assign regs_187_clock = clock; // @[:@130490.4]
  assign regs_187_reset = io_reset; // @[:@130491.4 RegFile.scala 76:16:@130498.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@130497.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@130501.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@130495.4]
  assign regs_188_clock = clock; // @[:@130504.4]
  assign regs_188_reset = io_reset; // @[:@130505.4 RegFile.scala 76:16:@130512.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@130511.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@130515.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@130509.4]
  assign regs_189_clock = clock; // @[:@130518.4]
  assign regs_189_reset = io_reset; // @[:@130519.4 RegFile.scala 76:16:@130526.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@130525.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@130529.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@130523.4]
  assign regs_190_clock = clock; // @[:@130532.4]
  assign regs_190_reset = io_reset; // @[:@130533.4 RegFile.scala 76:16:@130540.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@130539.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@130543.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@130537.4]
  assign regs_191_clock = clock; // @[:@130546.4]
  assign regs_191_reset = io_reset; // @[:@130547.4 RegFile.scala 76:16:@130554.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@130553.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@130557.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@130551.4]
  assign regs_192_clock = clock; // @[:@130560.4]
  assign regs_192_reset = io_reset; // @[:@130561.4 RegFile.scala 76:16:@130568.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@130567.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@130571.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@130565.4]
  assign regs_193_clock = clock; // @[:@130574.4]
  assign regs_193_reset = io_reset; // @[:@130575.4 RegFile.scala 76:16:@130582.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@130581.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@130585.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@130579.4]
  assign regs_194_clock = clock; // @[:@130588.4]
  assign regs_194_reset = io_reset; // @[:@130589.4 RegFile.scala 76:16:@130596.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@130595.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@130599.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@130593.4]
  assign regs_195_clock = clock; // @[:@130602.4]
  assign regs_195_reset = io_reset; // @[:@130603.4 RegFile.scala 76:16:@130610.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@130609.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@130613.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@130607.4]
  assign regs_196_clock = clock; // @[:@130616.4]
  assign regs_196_reset = io_reset; // @[:@130617.4 RegFile.scala 76:16:@130624.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@130623.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@130627.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@130621.4]
  assign regs_197_clock = clock; // @[:@130630.4]
  assign regs_197_reset = io_reset; // @[:@130631.4 RegFile.scala 76:16:@130638.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@130637.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@130641.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@130635.4]
  assign regs_198_clock = clock; // @[:@130644.4]
  assign regs_198_reset = io_reset; // @[:@130645.4 RegFile.scala 76:16:@130652.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@130651.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@130655.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@130649.4]
  assign regs_199_clock = clock; // @[:@130658.4]
  assign regs_199_reset = io_reset; // @[:@130659.4 RegFile.scala 76:16:@130666.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@130665.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@130669.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@130663.4]
  assign regs_200_clock = clock; // @[:@130672.4]
  assign regs_200_reset = io_reset; // @[:@130673.4 RegFile.scala 76:16:@130680.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@130679.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@130683.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@130677.4]
  assign regs_201_clock = clock; // @[:@130686.4]
  assign regs_201_reset = io_reset; // @[:@130687.4 RegFile.scala 76:16:@130694.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@130693.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@130697.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@130691.4]
  assign regs_202_clock = clock; // @[:@130700.4]
  assign regs_202_reset = io_reset; // @[:@130701.4 RegFile.scala 76:16:@130708.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@130707.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@130711.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@130705.4]
  assign regs_203_clock = clock; // @[:@130714.4]
  assign regs_203_reset = io_reset; // @[:@130715.4 RegFile.scala 76:16:@130722.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@130721.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@130725.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@130719.4]
  assign regs_204_clock = clock; // @[:@130728.4]
  assign regs_204_reset = io_reset; // @[:@130729.4 RegFile.scala 76:16:@130736.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@130735.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@130739.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@130733.4]
  assign regs_205_clock = clock; // @[:@130742.4]
  assign regs_205_reset = io_reset; // @[:@130743.4 RegFile.scala 76:16:@130750.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@130749.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@130753.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@130747.4]
  assign regs_206_clock = clock; // @[:@130756.4]
  assign regs_206_reset = io_reset; // @[:@130757.4 RegFile.scala 76:16:@130764.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@130763.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@130767.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@130761.4]
  assign regs_207_clock = clock; // @[:@130770.4]
  assign regs_207_reset = io_reset; // @[:@130771.4 RegFile.scala 76:16:@130778.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@130777.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@130781.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@130775.4]
  assign regs_208_clock = clock; // @[:@130784.4]
  assign regs_208_reset = io_reset; // @[:@130785.4 RegFile.scala 76:16:@130792.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@130791.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@130795.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@130789.4]
  assign regs_209_clock = clock; // @[:@130798.4]
  assign regs_209_reset = io_reset; // @[:@130799.4 RegFile.scala 76:16:@130806.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@130805.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@130809.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@130803.4]
  assign regs_210_clock = clock; // @[:@130812.4]
  assign regs_210_reset = io_reset; // @[:@130813.4 RegFile.scala 76:16:@130820.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@130819.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@130823.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@130817.4]
  assign regs_211_clock = clock; // @[:@130826.4]
  assign regs_211_reset = io_reset; // @[:@130827.4 RegFile.scala 76:16:@130834.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@130833.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@130837.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@130831.4]
  assign regs_212_clock = clock; // @[:@130840.4]
  assign regs_212_reset = io_reset; // @[:@130841.4 RegFile.scala 76:16:@130848.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@130847.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@130851.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@130845.4]
  assign regs_213_clock = clock; // @[:@130854.4]
  assign regs_213_reset = io_reset; // @[:@130855.4 RegFile.scala 76:16:@130862.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@130861.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@130865.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@130859.4]
  assign regs_214_clock = clock; // @[:@130868.4]
  assign regs_214_reset = io_reset; // @[:@130869.4 RegFile.scala 76:16:@130876.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@130875.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@130879.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@130873.4]
  assign regs_215_clock = clock; // @[:@130882.4]
  assign regs_215_reset = io_reset; // @[:@130883.4 RegFile.scala 76:16:@130890.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@130889.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@130893.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@130887.4]
  assign regs_216_clock = clock; // @[:@130896.4]
  assign regs_216_reset = io_reset; // @[:@130897.4 RegFile.scala 76:16:@130904.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@130903.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@130907.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@130901.4]
  assign regs_217_clock = clock; // @[:@130910.4]
  assign regs_217_reset = io_reset; // @[:@130911.4 RegFile.scala 76:16:@130918.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@130917.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@130921.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@130915.4]
  assign regs_218_clock = clock; // @[:@130924.4]
  assign regs_218_reset = io_reset; // @[:@130925.4 RegFile.scala 76:16:@130932.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@130931.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@130935.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@130929.4]
  assign regs_219_clock = clock; // @[:@130938.4]
  assign regs_219_reset = io_reset; // @[:@130939.4 RegFile.scala 76:16:@130946.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@130945.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@130949.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@130943.4]
  assign regs_220_clock = clock; // @[:@130952.4]
  assign regs_220_reset = io_reset; // @[:@130953.4 RegFile.scala 76:16:@130960.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@130959.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@130963.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@130957.4]
  assign regs_221_clock = clock; // @[:@130966.4]
  assign regs_221_reset = io_reset; // @[:@130967.4 RegFile.scala 76:16:@130974.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@130973.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@130977.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@130971.4]
  assign regs_222_clock = clock; // @[:@130980.4]
  assign regs_222_reset = io_reset; // @[:@130981.4 RegFile.scala 76:16:@130988.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@130987.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@130991.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@130985.4]
  assign regs_223_clock = clock; // @[:@130994.4]
  assign regs_223_reset = io_reset; // @[:@130995.4 RegFile.scala 76:16:@131002.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@131001.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@131005.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@130999.4]
  assign regs_224_clock = clock; // @[:@131008.4]
  assign regs_224_reset = io_reset; // @[:@131009.4 RegFile.scala 76:16:@131016.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@131015.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@131019.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@131013.4]
  assign regs_225_clock = clock; // @[:@131022.4]
  assign regs_225_reset = io_reset; // @[:@131023.4 RegFile.scala 76:16:@131030.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@131029.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@131033.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@131027.4]
  assign regs_226_clock = clock; // @[:@131036.4]
  assign regs_226_reset = io_reset; // @[:@131037.4 RegFile.scala 76:16:@131044.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@131043.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@131047.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@131041.4]
  assign regs_227_clock = clock; // @[:@131050.4]
  assign regs_227_reset = io_reset; // @[:@131051.4 RegFile.scala 76:16:@131058.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@131057.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@131061.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@131055.4]
  assign regs_228_clock = clock; // @[:@131064.4]
  assign regs_228_reset = io_reset; // @[:@131065.4 RegFile.scala 76:16:@131072.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@131071.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@131075.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@131069.4]
  assign regs_229_clock = clock; // @[:@131078.4]
  assign regs_229_reset = io_reset; // @[:@131079.4 RegFile.scala 76:16:@131086.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@131085.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@131089.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@131083.4]
  assign regs_230_clock = clock; // @[:@131092.4]
  assign regs_230_reset = io_reset; // @[:@131093.4 RegFile.scala 76:16:@131100.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@131099.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@131103.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@131097.4]
  assign regs_231_clock = clock; // @[:@131106.4]
  assign regs_231_reset = io_reset; // @[:@131107.4 RegFile.scala 76:16:@131114.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@131113.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@131117.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@131111.4]
  assign regs_232_clock = clock; // @[:@131120.4]
  assign regs_232_reset = io_reset; // @[:@131121.4 RegFile.scala 76:16:@131128.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@131127.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@131131.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@131125.4]
  assign regs_233_clock = clock; // @[:@131134.4]
  assign regs_233_reset = io_reset; // @[:@131135.4 RegFile.scala 76:16:@131142.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@131141.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@131145.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@131139.4]
  assign regs_234_clock = clock; // @[:@131148.4]
  assign regs_234_reset = io_reset; // @[:@131149.4 RegFile.scala 76:16:@131156.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@131155.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@131159.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@131153.4]
  assign regs_235_clock = clock; // @[:@131162.4]
  assign regs_235_reset = io_reset; // @[:@131163.4 RegFile.scala 76:16:@131170.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@131169.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@131173.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@131167.4]
  assign regs_236_clock = clock; // @[:@131176.4]
  assign regs_236_reset = io_reset; // @[:@131177.4 RegFile.scala 76:16:@131184.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@131183.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@131187.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@131181.4]
  assign regs_237_clock = clock; // @[:@131190.4]
  assign regs_237_reset = io_reset; // @[:@131191.4 RegFile.scala 76:16:@131198.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@131197.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@131201.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@131195.4]
  assign regs_238_clock = clock; // @[:@131204.4]
  assign regs_238_reset = io_reset; // @[:@131205.4 RegFile.scala 76:16:@131212.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@131211.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@131215.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@131209.4]
  assign regs_239_clock = clock; // @[:@131218.4]
  assign regs_239_reset = io_reset; // @[:@131219.4 RegFile.scala 76:16:@131226.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@131225.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@131229.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@131223.4]
  assign regs_240_clock = clock; // @[:@131232.4]
  assign regs_240_reset = io_reset; // @[:@131233.4 RegFile.scala 76:16:@131240.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@131239.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@131243.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@131237.4]
  assign regs_241_clock = clock; // @[:@131246.4]
  assign regs_241_reset = io_reset; // @[:@131247.4 RegFile.scala 76:16:@131254.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@131253.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@131257.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@131251.4]
  assign regs_242_clock = clock; // @[:@131260.4]
  assign regs_242_reset = io_reset; // @[:@131261.4 RegFile.scala 76:16:@131268.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@131267.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@131271.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@131265.4]
  assign regs_243_clock = clock; // @[:@131274.4]
  assign regs_243_reset = io_reset; // @[:@131275.4 RegFile.scala 76:16:@131282.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@131281.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@131285.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@131279.4]
  assign regs_244_clock = clock; // @[:@131288.4]
  assign regs_244_reset = io_reset; // @[:@131289.4 RegFile.scala 76:16:@131296.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@131295.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@131299.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@131293.4]
  assign regs_245_clock = clock; // @[:@131302.4]
  assign regs_245_reset = io_reset; // @[:@131303.4 RegFile.scala 76:16:@131310.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@131309.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@131313.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@131307.4]
  assign regs_246_clock = clock; // @[:@131316.4]
  assign regs_246_reset = io_reset; // @[:@131317.4 RegFile.scala 76:16:@131324.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@131323.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@131327.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@131321.4]
  assign regs_247_clock = clock; // @[:@131330.4]
  assign regs_247_reset = io_reset; // @[:@131331.4 RegFile.scala 76:16:@131338.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@131337.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@131341.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@131335.4]
  assign regs_248_clock = clock; // @[:@131344.4]
  assign regs_248_reset = io_reset; // @[:@131345.4 RegFile.scala 76:16:@131352.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@131351.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@131355.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@131349.4]
  assign regs_249_clock = clock; // @[:@131358.4]
  assign regs_249_reset = io_reset; // @[:@131359.4 RegFile.scala 76:16:@131366.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@131365.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@131369.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@131363.4]
  assign regs_250_clock = clock; // @[:@131372.4]
  assign regs_250_reset = io_reset; // @[:@131373.4 RegFile.scala 76:16:@131380.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@131379.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@131383.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@131377.4]
  assign regs_251_clock = clock; // @[:@131386.4]
  assign regs_251_reset = io_reset; // @[:@131387.4 RegFile.scala 76:16:@131394.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@131393.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@131397.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@131391.4]
  assign regs_252_clock = clock; // @[:@131400.4]
  assign regs_252_reset = io_reset; // @[:@131401.4 RegFile.scala 76:16:@131408.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@131407.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@131411.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@131405.4]
  assign regs_253_clock = clock; // @[:@131414.4]
  assign regs_253_reset = io_reset; // @[:@131415.4 RegFile.scala 76:16:@131422.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@131421.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@131425.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@131419.4]
  assign regs_254_clock = clock; // @[:@131428.4]
  assign regs_254_reset = io_reset; // @[:@131429.4 RegFile.scala 76:16:@131436.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@131435.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@131439.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@131433.4]
  assign regs_255_clock = clock; // @[:@131442.4]
  assign regs_255_reset = io_reset; // @[:@131443.4 RegFile.scala 76:16:@131450.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@131449.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@131453.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@131447.4]
  assign regs_256_clock = clock; // @[:@131456.4]
  assign regs_256_reset = io_reset; // @[:@131457.4 RegFile.scala 76:16:@131464.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@131463.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@131467.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@131461.4]
  assign regs_257_clock = clock; // @[:@131470.4]
  assign regs_257_reset = io_reset; // @[:@131471.4 RegFile.scala 76:16:@131478.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@131477.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@131481.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@131475.4]
  assign regs_258_clock = clock; // @[:@131484.4]
  assign regs_258_reset = io_reset; // @[:@131485.4 RegFile.scala 76:16:@131492.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@131491.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@131495.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@131489.4]
  assign regs_259_clock = clock; // @[:@131498.4]
  assign regs_259_reset = io_reset; // @[:@131499.4 RegFile.scala 76:16:@131506.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@131505.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@131509.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@131503.4]
  assign regs_260_clock = clock; // @[:@131512.4]
  assign regs_260_reset = io_reset; // @[:@131513.4 RegFile.scala 76:16:@131520.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@131519.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@131523.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@131517.4]
  assign regs_261_clock = clock; // @[:@131526.4]
  assign regs_261_reset = io_reset; // @[:@131527.4 RegFile.scala 76:16:@131534.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@131533.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@131537.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@131531.4]
  assign regs_262_clock = clock; // @[:@131540.4]
  assign regs_262_reset = io_reset; // @[:@131541.4 RegFile.scala 76:16:@131548.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@131547.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@131551.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@131545.4]
  assign regs_263_clock = clock; // @[:@131554.4]
  assign regs_263_reset = io_reset; // @[:@131555.4 RegFile.scala 76:16:@131562.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@131561.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@131565.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@131559.4]
  assign regs_264_clock = clock; // @[:@131568.4]
  assign regs_264_reset = io_reset; // @[:@131569.4 RegFile.scala 76:16:@131576.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@131575.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@131579.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@131573.4]
  assign regs_265_clock = clock; // @[:@131582.4]
  assign regs_265_reset = io_reset; // @[:@131583.4 RegFile.scala 76:16:@131590.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@131589.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@131593.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@131587.4]
  assign regs_266_clock = clock; // @[:@131596.4]
  assign regs_266_reset = io_reset; // @[:@131597.4 RegFile.scala 76:16:@131604.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@131603.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@131607.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@131601.4]
  assign regs_267_clock = clock; // @[:@131610.4]
  assign regs_267_reset = io_reset; // @[:@131611.4 RegFile.scala 76:16:@131618.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@131617.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@131621.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@131615.4]
  assign regs_268_clock = clock; // @[:@131624.4]
  assign regs_268_reset = io_reset; // @[:@131625.4 RegFile.scala 76:16:@131632.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@131631.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@131635.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@131629.4]
  assign regs_269_clock = clock; // @[:@131638.4]
  assign regs_269_reset = io_reset; // @[:@131639.4 RegFile.scala 76:16:@131646.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@131645.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@131649.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@131643.4]
  assign regs_270_clock = clock; // @[:@131652.4]
  assign regs_270_reset = io_reset; // @[:@131653.4 RegFile.scala 76:16:@131660.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@131659.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@131663.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@131657.4]
  assign regs_271_clock = clock; // @[:@131666.4]
  assign regs_271_reset = io_reset; // @[:@131667.4 RegFile.scala 76:16:@131674.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@131673.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@131677.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@131671.4]
  assign regs_272_clock = clock; // @[:@131680.4]
  assign regs_272_reset = io_reset; // @[:@131681.4 RegFile.scala 76:16:@131688.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@131687.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@131691.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@131685.4]
  assign regs_273_clock = clock; // @[:@131694.4]
  assign regs_273_reset = io_reset; // @[:@131695.4 RegFile.scala 76:16:@131702.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@131701.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@131705.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@131699.4]
  assign regs_274_clock = clock; // @[:@131708.4]
  assign regs_274_reset = io_reset; // @[:@131709.4 RegFile.scala 76:16:@131716.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@131715.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@131719.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@131713.4]
  assign regs_275_clock = clock; // @[:@131722.4]
  assign regs_275_reset = io_reset; // @[:@131723.4 RegFile.scala 76:16:@131730.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@131729.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@131733.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@131727.4]
  assign regs_276_clock = clock; // @[:@131736.4]
  assign regs_276_reset = io_reset; // @[:@131737.4 RegFile.scala 76:16:@131744.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@131743.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@131747.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@131741.4]
  assign regs_277_clock = clock; // @[:@131750.4]
  assign regs_277_reset = io_reset; // @[:@131751.4 RegFile.scala 76:16:@131758.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@131757.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@131761.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@131755.4]
  assign regs_278_clock = clock; // @[:@131764.4]
  assign regs_278_reset = io_reset; // @[:@131765.4 RegFile.scala 76:16:@131772.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@131771.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@131775.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@131769.4]
  assign regs_279_clock = clock; // @[:@131778.4]
  assign regs_279_reset = io_reset; // @[:@131779.4 RegFile.scala 76:16:@131786.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@131785.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@131789.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@131783.4]
  assign regs_280_clock = clock; // @[:@131792.4]
  assign regs_280_reset = io_reset; // @[:@131793.4 RegFile.scala 76:16:@131800.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@131799.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@131803.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@131797.4]
  assign regs_281_clock = clock; // @[:@131806.4]
  assign regs_281_reset = io_reset; // @[:@131807.4 RegFile.scala 76:16:@131814.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@131813.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@131817.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@131811.4]
  assign regs_282_clock = clock; // @[:@131820.4]
  assign regs_282_reset = io_reset; // @[:@131821.4 RegFile.scala 76:16:@131828.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@131827.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@131831.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@131825.4]
  assign regs_283_clock = clock; // @[:@131834.4]
  assign regs_283_reset = io_reset; // @[:@131835.4 RegFile.scala 76:16:@131842.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@131841.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@131845.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@131839.4]
  assign regs_284_clock = clock; // @[:@131848.4]
  assign regs_284_reset = io_reset; // @[:@131849.4 RegFile.scala 76:16:@131856.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@131855.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@131859.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@131853.4]
  assign regs_285_clock = clock; // @[:@131862.4]
  assign regs_285_reset = io_reset; // @[:@131863.4 RegFile.scala 76:16:@131870.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@131869.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@131873.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@131867.4]
  assign regs_286_clock = clock; // @[:@131876.4]
  assign regs_286_reset = io_reset; // @[:@131877.4 RegFile.scala 76:16:@131884.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@131883.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@131887.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@131881.4]
  assign regs_287_clock = clock; // @[:@131890.4]
  assign regs_287_reset = io_reset; // @[:@131891.4 RegFile.scala 76:16:@131898.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@131897.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@131901.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@131895.4]
  assign regs_288_clock = clock; // @[:@131904.4]
  assign regs_288_reset = io_reset; // @[:@131905.4 RegFile.scala 76:16:@131912.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@131911.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@131915.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@131909.4]
  assign regs_289_clock = clock; // @[:@131918.4]
  assign regs_289_reset = io_reset; // @[:@131919.4 RegFile.scala 76:16:@131926.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@131925.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@131929.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@131923.4]
  assign regs_290_clock = clock; // @[:@131932.4]
  assign regs_290_reset = io_reset; // @[:@131933.4 RegFile.scala 76:16:@131940.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@131939.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@131943.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@131937.4]
  assign regs_291_clock = clock; // @[:@131946.4]
  assign regs_291_reset = io_reset; // @[:@131947.4 RegFile.scala 76:16:@131954.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@131953.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@131957.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@131951.4]
  assign regs_292_clock = clock; // @[:@131960.4]
  assign regs_292_reset = io_reset; // @[:@131961.4 RegFile.scala 76:16:@131968.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@131967.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@131971.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@131965.4]
  assign regs_293_clock = clock; // @[:@131974.4]
  assign regs_293_reset = io_reset; // @[:@131975.4 RegFile.scala 76:16:@131982.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@131981.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@131985.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@131979.4]
  assign regs_294_clock = clock; // @[:@131988.4]
  assign regs_294_reset = io_reset; // @[:@131989.4 RegFile.scala 76:16:@131996.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@131995.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@131999.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@131993.4]
  assign regs_295_clock = clock; // @[:@132002.4]
  assign regs_295_reset = io_reset; // @[:@132003.4 RegFile.scala 76:16:@132010.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@132009.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@132013.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@132007.4]
  assign regs_296_clock = clock; // @[:@132016.4]
  assign regs_296_reset = io_reset; // @[:@132017.4 RegFile.scala 76:16:@132024.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@132023.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@132027.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@132021.4]
  assign regs_297_clock = clock; // @[:@132030.4]
  assign regs_297_reset = io_reset; // @[:@132031.4 RegFile.scala 76:16:@132038.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@132037.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@132041.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@132035.4]
  assign regs_298_clock = clock; // @[:@132044.4]
  assign regs_298_reset = io_reset; // @[:@132045.4 RegFile.scala 76:16:@132052.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@132051.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@132055.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@132049.4]
  assign regs_299_clock = clock; // @[:@132058.4]
  assign regs_299_reset = io_reset; // @[:@132059.4 RegFile.scala 76:16:@132066.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@132065.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@132069.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@132063.4]
  assign regs_300_clock = clock; // @[:@132072.4]
  assign regs_300_reset = io_reset; // @[:@132073.4 RegFile.scala 76:16:@132080.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@132079.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@132083.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@132077.4]
  assign regs_301_clock = clock; // @[:@132086.4]
  assign regs_301_reset = io_reset; // @[:@132087.4 RegFile.scala 76:16:@132094.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@132093.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@132097.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@132091.4]
  assign regs_302_clock = clock; // @[:@132100.4]
  assign regs_302_reset = io_reset; // @[:@132101.4 RegFile.scala 76:16:@132108.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@132107.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@132111.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@132105.4]
  assign regs_303_clock = clock; // @[:@132114.4]
  assign regs_303_reset = io_reset; // @[:@132115.4 RegFile.scala 76:16:@132122.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@132121.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@132125.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@132119.4]
  assign regs_304_clock = clock; // @[:@132128.4]
  assign regs_304_reset = io_reset; // @[:@132129.4 RegFile.scala 76:16:@132136.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@132135.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@132139.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@132133.4]
  assign regs_305_clock = clock; // @[:@132142.4]
  assign regs_305_reset = io_reset; // @[:@132143.4 RegFile.scala 76:16:@132150.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@132149.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@132153.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@132147.4]
  assign regs_306_clock = clock; // @[:@132156.4]
  assign regs_306_reset = io_reset; // @[:@132157.4 RegFile.scala 76:16:@132164.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@132163.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@132167.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@132161.4]
  assign regs_307_clock = clock; // @[:@132170.4]
  assign regs_307_reset = io_reset; // @[:@132171.4 RegFile.scala 76:16:@132178.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@132177.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@132181.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@132175.4]
  assign regs_308_clock = clock; // @[:@132184.4]
  assign regs_308_reset = io_reset; // @[:@132185.4 RegFile.scala 76:16:@132192.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@132191.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@132195.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@132189.4]
  assign regs_309_clock = clock; // @[:@132198.4]
  assign regs_309_reset = io_reset; // @[:@132199.4 RegFile.scala 76:16:@132206.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@132205.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@132209.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@132203.4]
  assign regs_310_clock = clock; // @[:@132212.4]
  assign regs_310_reset = io_reset; // @[:@132213.4 RegFile.scala 76:16:@132220.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@132219.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@132223.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@132217.4]
  assign regs_311_clock = clock; // @[:@132226.4]
  assign regs_311_reset = io_reset; // @[:@132227.4 RegFile.scala 76:16:@132234.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@132233.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@132237.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@132231.4]
  assign regs_312_clock = clock; // @[:@132240.4]
  assign regs_312_reset = io_reset; // @[:@132241.4 RegFile.scala 76:16:@132248.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@132247.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@132251.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@132245.4]
  assign regs_313_clock = clock; // @[:@132254.4]
  assign regs_313_reset = io_reset; // @[:@132255.4 RegFile.scala 76:16:@132262.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@132261.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@132265.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@132259.4]
  assign regs_314_clock = clock; // @[:@132268.4]
  assign regs_314_reset = io_reset; // @[:@132269.4 RegFile.scala 76:16:@132276.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@132275.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@132279.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@132273.4]
  assign regs_315_clock = clock; // @[:@132282.4]
  assign regs_315_reset = io_reset; // @[:@132283.4 RegFile.scala 76:16:@132290.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@132289.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@132293.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@132287.4]
  assign regs_316_clock = clock; // @[:@132296.4]
  assign regs_316_reset = io_reset; // @[:@132297.4 RegFile.scala 76:16:@132304.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@132303.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@132307.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@132301.4]
  assign regs_317_clock = clock; // @[:@132310.4]
  assign regs_317_reset = io_reset; // @[:@132311.4 RegFile.scala 76:16:@132318.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@132317.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@132321.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@132315.4]
  assign regs_318_clock = clock; // @[:@132324.4]
  assign regs_318_reset = io_reset; // @[:@132325.4 RegFile.scala 76:16:@132332.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@132331.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@132335.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@132329.4]
  assign regs_319_clock = clock; // @[:@132338.4]
  assign regs_319_reset = io_reset; // @[:@132339.4 RegFile.scala 76:16:@132346.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@132345.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@132349.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@132343.4]
  assign regs_320_clock = clock; // @[:@132352.4]
  assign regs_320_reset = io_reset; // @[:@132353.4 RegFile.scala 76:16:@132360.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@132359.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@132363.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@132357.4]
  assign regs_321_clock = clock; // @[:@132366.4]
  assign regs_321_reset = io_reset; // @[:@132367.4 RegFile.scala 76:16:@132374.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@132373.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@132377.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@132371.4]
  assign regs_322_clock = clock; // @[:@132380.4]
  assign regs_322_reset = io_reset; // @[:@132381.4 RegFile.scala 76:16:@132388.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@132387.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@132391.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@132385.4]
  assign regs_323_clock = clock; // @[:@132394.4]
  assign regs_323_reset = io_reset; // @[:@132395.4 RegFile.scala 76:16:@132402.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@132401.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@132405.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@132399.4]
  assign regs_324_clock = clock; // @[:@132408.4]
  assign regs_324_reset = io_reset; // @[:@132409.4 RegFile.scala 76:16:@132416.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@132415.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@132419.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@132413.4]
  assign regs_325_clock = clock; // @[:@132422.4]
  assign regs_325_reset = io_reset; // @[:@132423.4 RegFile.scala 76:16:@132430.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@132429.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@132433.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@132427.4]
  assign regs_326_clock = clock; // @[:@132436.4]
  assign regs_326_reset = io_reset; // @[:@132437.4 RegFile.scala 76:16:@132444.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@132443.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@132447.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@132441.4]
  assign regs_327_clock = clock; // @[:@132450.4]
  assign regs_327_reset = io_reset; // @[:@132451.4 RegFile.scala 76:16:@132458.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@132457.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@132461.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@132455.4]
  assign regs_328_clock = clock; // @[:@132464.4]
  assign regs_328_reset = io_reset; // @[:@132465.4 RegFile.scala 76:16:@132472.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@132471.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@132475.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@132469.4]
  assign regs_329_clock = clock; // @[:@132478.4]
  assign regs_329_reset = io_reset; // @[:@132479.4 RegFile.scala 76:16:@132486.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@132485.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@132489.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@132483.4]
  assign regs_330_clock = clock; // @[:@132492.4]
  assign regs_330_reset = io_reset; // @[:@132493.4 RegFile.scala 76:16:@132500.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@132499.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@132503.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@132497.4]
  assign regs_331_clock = clock; // @[:@132506.4]
  assign regs_331_reset = io_reset; // @[:@132507.4 RegFile.scala 76:16:@132514.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@132513.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@132517.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@132511.4]
  assign regs_332_clock = clock; // @[:@132520.4]
  assign regs_332_reset = io_reset; // @[:@132521.4 RegFile.scala 76:16:@132528.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@132527.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@132531.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@132525.4]
  assign regs_333_clock = clock; // @[:@132534.4]
  assign regs_333_reset = io_reset; // @[:@132535.4 RegFile.scala 76:16:@132542.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@132541.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@132545.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@132539.4]
  assign regs_334_clock = clock; // @[:@132548.4]
  assign regs_334_reset = io_reset; // @[:@132549.4 RegFile.scala 76:16:@132556.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@132555.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@132559.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@132553.4]
  assign regs_335_clock = clock; // @[:@132562.4]
  assign regs_335_reset = io_reset; // @[:@132563.4 RegFile.scala 76:16:@132570.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@132569.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@132573.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@132567.4]
  assign regs_336_clock = clock; // @[:@132576.4]
  assign regs_336_reset = io_reset; // @[:@132577.4 RegFile.scala 76:16:@132584.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@132583.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@132587.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@132581.4]
  assign regs_337_clock = clock; // @[:@132590.4]
  assign regs_337_reset = io_reset; // @[:@132591.4 RegFile.scala 76:16:@132598.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@132597.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@132601.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@132595.4]
  assign regs_338_clock = clock; // @[:@132604.4]
  assign regs_338_reset = io_reset; // @[:@132605.4 RegFile.scala 76:16:@132612.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@132611.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@132615.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@132609.4]
  assign regs_339_clock = clock; // @[:@132618.4]
  assign regs_339_reset = io_reset; // @[:@132619.4 RegFile.scala 76:16:@132626.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@132625.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@132629.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@132623.4]
  assign regs_340_clock = clock; // @[:@132632.4]
  assign regs_340_reset = io_reset; // @[:@132633.4 RegFile.scala 76:16:@132640.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@132639.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@132643.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@132637.4]
  assign regs_341_clock = clock; // @[:@132646.4]
  assign regs_341_reset = io_reset; // @[:@132647.4 RegFile.scala 76:16:@132654.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@132653.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@132657.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@132651.4]
  assign regs_342_clock = clock; // @[:@132660.4]
  assign regs_342_reset = io_reset; // @[:@132661.4 RegFile.scala 76:16:@132668.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@132667.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@132671.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@132665.4]
  assign regs_343_clock = clock; // @[:@132674.4]
  assign regs_343_reset = io_reset; // @[:@132675.4 RegFile.scala 76:16:@132682.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@132681.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@132685.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@132679.4]
  assign regs_344_clock = clock; // @[:@132688.4]
  assign regs_344_reset = io_reset; // @[:@132689.4 RegFile.scala 76:16:@132696.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@132695.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@132699.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@132693.4]
  assign regs_345_clock = clock; // @[:@132702.4]
  assign regs_345_reset = io_reset; // @[:@132703.4 RegFile.scala 76:16:@132710.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@132709.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@132713.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@132707.4]
  assign regs_346_clock = clock; // @[:@132716.4]
  assign regs_346_reset = io_reset; // @[:@132717.4 RegFile.scala 76:16:@132724.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@132723.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@132727.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@132721.4]
  assign regs_347_clock = clock; // @[:@132730.4]
  assign regs_347_reset = io_reset; // @[:@132731.4 RegFile.scala 76:16:@132738.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@132737.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@132741.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@132735.4]
  assign regs_348_clock = clock; // @[:@132744.4]
  assign regs_348_reset = io_reset; // @[:@132745.4 RegFile.scala 76:16:@132752.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@132751.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@132755.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@132749.4]
  assign regs_349_clock = clock; // @[:@132758.4]
  assign regs_349_reset = io_reset; // @[:@132759.4 RegFile.scala 76:16:@132766.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@132765.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@132769.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@132763.4]
  assign regs_350_clock = clock; // @[:@132772.4]
  assign regs_350_reset = io_reset; // @[:@132773.4 RegFile.scala 76:16:@132780.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@132779.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@132783.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@132777.4]
  assign regs_351_clock = clock; // @[:@132786.4]
  assign regs_351_reset = io_reset; // @[:@132787.4 RegFile.scala 76:16:@132794.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@132793.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@132797.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@132791.4]
  assign regs_352_clock = clock; // @[:@132800.4]
  assign regs_352_reset = io_reset; // @[:@132801.4 RegFile.scala 76:16:@132808.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@132807.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@132811.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@132805.4]
  assign regs_353_clock = clock; // @[:@132814.4]
  assign regs_353_reset = io_reset; // @[:@132815.4 RegFile.scala 76:16:@132822.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@132821.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@132825.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@132819.4]
  assign regs_354_clock = clock; // @[:@132828.4]
  assign regs_354_reset = io_reset; // @[:@132829.4 RegFile.scala 76:16:@132836.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@132835.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@132839.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@132833.4]
  assign regs_355_clock = clock; // @[:@132842.4]
  assign regs_355_reset = io_reset; // @[:@132843.4 RegFile.scala 76:16:@132850.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@132849.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@132853.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@132847.4]
  assign regs_356_clock = clock; // @[:@132856.4]
  assign regs_356_reset = io_reset; // @[:@132857.4 RegFile.scala 76:16:@132864.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@132863.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@132867.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@132861.4]
  assign regs_357_clock = clock; // @[:@132870.4]
  assign regs_357_reset = io_reset; // @[:@132871.4 RegFile.scala 76:16:@132878.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@132877.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@132881.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@132875.4]
  assign regs_358_clock = clock; // @[:@132884.4]
  assign regs_358_reset = io_reset; // @[:@132885.4 RegFile.scala 76:16:@132892.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@132891.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@132895.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@132889.4]
  assign regs_359_clock = clock; // @[:@132898.4]
  assign regs_359_reset = io_reset; // @[:@132899.4 RegFile.scala 76:16:@132906.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@132905.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@132909.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@132903.4]
  assign regs_360_clock = clock; // @[:@132912.4]
  assign regs_360_reset = io_reset; // @[:@132913.4 RegFile.scala 76:16:@132920.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@132919.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@132923.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@132917.4]
  assign regs_361_clock = clock; // @[:@132926.4]
  assign regs_361_reset = io_reset; // @[:@132927.4 RegFile.scala 76:16:@132934.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@132933.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@132937.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@132931.4]
  assign regs_362_clock = clock; // @[:@132940.4]
  assign regs_362_reset = io_reset; // @[:@132941.4 RegFile.scala 76:16:@132948.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@132947.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@132951.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@132945.4]
  assign regs_363_clock = clock; // @[:@132954.4]
  assign regs_363_reset = io_reset; // @[:@132955.4 RegFile.scala 76:16:@132962.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@132961.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@132965.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@132959.4]
  assign regs_364_clock = clock; // @[:@132968.4]
  assign regs_364_reset = io_reset; // @[:@132969.4 RegFile.scala 76:16:@132976.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@132975.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@132979.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@132973.4]
  assign regs_365_clock = clock; // @[:@132982.4]
  assign regs_365_reset = io_reset; // @[:@132983.4 RegFile.scala 76:16:@132990.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@132989.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@132993.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@132987.4]
  assign regs_366_clock = clock; // @[:@132996.4]
  assign regs_366_reset = io_reset; // @[:@132997.4 RegFile.scala 76:16:@133004.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@133003.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@133007.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@133001.4]
  assign regs_367_clock = clock; // @[:@133010.4]
  assign regs_367_reset = io_reset; // @[:@133011.4 RegFile.scala 76:16:@133018.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@133017.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@133021.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@133015.4]
  assign regs_368_clock = clock; // @[:@133024.4]
  assign regs_368_reset = io_reset; // @[:@133025.4 RegFile.scala 76:16:@133032.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@133031.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@133035.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@133029.4]
  assign regs_369_clock = clock; // @[:@133038.4]
  assign regs_369_reset = io_reset; // @[:@133039.4 RegFile.scala 76:16:@133046.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@133045.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@133049.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@133043.4]
  assign regs_370_clock = clock; // @[:@133052.4]
  assign regs_370_reset = io_reset; // @[:@133053.4 RegFile.scala 76:16:@133060.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@133059.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@133063.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@133057.4]
  assign regs_371_clock = clock; // @[:@133066.4]
  assign regs_371_reset = io_reset; // @[:@133067.4 RegFile.scala 76:16:@133074.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@133073.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@133077.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@133071.4]
  assign regs_372_clock = clock; // @[:@133080.4]
  assign regs_372_reset = io_reset; // @[:@133081.4 RegFile.scala 76:16:@133088.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@133087.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@133091.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@133085.4]
  assign regs_373_clock = clock; // @[:@133094.4]
  assign regs_373_reset = io_reset; // @[:@133095.4 RegFile.scala 76:16:@133102.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@133101.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@133105.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@133099.4]
  assign regs_374_clock = clock; // @[:@133108.4]
  assign regs_374_reset = io_reset; // @[:@133109.4 RegFile.scala 76:16:@133116.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@133115.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@133119.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@133113.4]
  assign regs_375_clock = clock; // @[:@133122.4]
  assign regs_375_reset = io_reset; // @[:@133123.4 RegFile.scala 76:16:@133130.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@133129.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@133133.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@133127.4]
  assign regs_376_clock = clock; // @[:@133136.4]
  assign regs_376_reset = io_reset; // @[:@133137.4 RegFile.scala 76:16:@133144.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@133143.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@133147.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@133141.4]
  assign regs_377_clock = clock; // @[:@133150.4]
  assign regs_377_reset = io_reset; // @[:@133151.4 RegFile.scala 76:16:@133158.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@133157.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@133161.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@133155.4]
  assign regs_378_clock = clock; // @[:@133164.4]
  assign regs_378_reset = io_reset; // @[:@133165.4 RegFile.scala 76:16:@133172.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@133171.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@133175.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@133169.4]
  assign regs_379_clock = clock; // @[:@133178.4]
  assign regs_379_reset = io_reset; // @[:@133179.4 RegFile.scala 76:16:@133186.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@133185.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@133189.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@133183.4]
  assign regs_380_clock = clock; // @[:@133192.4]
  assign regs_380_reset = io_reset; // @[:@133193.4 RegFile.scala 76:16:@133200.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@133199.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@133203.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@133197.4]
  assign regs_381_clock = clock; // @[:@133206.4]
  assign regs_381_reset = io_reset; // @[:@133207.4 RegFile.scala 76:16:@133214.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@133213.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@133217.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@133211.4]
  assign regs_382_clock = clock; // @[:@133220.4]
  assign regs_382_reset = io_reset; // @[:@133221.4 RegFile.scala 76:16:@133228.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@133227.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@133231.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@133225.4]
  assign regs_383_clock = clock; // @[:@133234.4]
  assign regs_383_reset = io_reset; // @[:@133235.4 RegFile.scala 76:16:@133242.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@133241.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@133245.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@133239.4]
  assign regs_384_clock = clock; // @[:@133248.4]
  assign regs_384_reset = io_reset; // @[:@133249.4 RegFile.scala 76:16:@133256.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@133255.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@133259.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@133253.4]
  assign regs_385_clock = clock; // @[:@133262.4]
  assign regs_385_reset = io_reset; // @[:@133263.4 RegFile.scala 76:16:@133270.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@133269.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@133273.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@133267.4]
  assign regs_386_clock = clock; // @[:@133276.4]
  assign regs_386_reset = io_reset; // @[:@133277.4 RegFile.scala 76:16:@133284.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@133283.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@133287.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@133281.4]
  assign regs_387_clock = clock; // @[:@133290.4]
  assign regs_387_reset = io_reset; // @[:@133291.4 RegFile.scala 76:16:@133298.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@133297.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@133301.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@133295.4]
  assign regs_388_clock = clock; // @[:@133304.4]
  assign regs_388_reset = io_reset; // @[:@133305.4 RegFile.scala 76:16:@133312.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@133311.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@133315.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@133309.4]
  assign regs_389_clock = clock; // @[:@133318.4]
  assign regs_389_reset = io_reset; // @[:@133319.4 RegFile.scala 76:16:@133326.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@133325.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@133329.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@133323.4]
  assign regs_390_clock = clock; // @[:@133332.4]
  assign regs_390_reset = io_reset; // @[:@133333.4 RegFile.scala 76:16:@133340.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@133339.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@133343.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@133337.4]
  assign regs_391_clock = clock; // @[:@133346.4]
  assign regs_391_reset = io_reset; // @[:@133347.4 RegFile.scala 76:16:@133354.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@133353.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@133357.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@133351.4]
  assign regs_392_clock = clock; // @[:@133360.4]
  assign regs_392_reset = io_reset; // @[:@133361.4 RegFile.scala 76:16:@133368.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@133367.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@133371.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@133365.4]
  assign regs_393_clock = clock; // @[:@133374.4]
  assign regs_393_reset = io_reset; // @[:@133375.4 RegFile.scala 76:16:@133382.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@133381.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@133385.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@133379.4]
  assign regs_394_clock = clock; // @[:@133388.4]
  assign regs_394_reset = io_reset; // @[:@133389.4 RegFile.scala 76:16:@133396.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@133395.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@133399.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@133393.4]
  assign regs_395_clock = clock; // @[:@133402.4]
  assign regs_395_reset = io_reset; // @[:@133403.4 RegFile.scala 76:16:@133410.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@133409.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@133413.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@133407.4]
  assign regs_396_clock = clock; // @[:@133416.4]
  assign regs_396_reset = io_reset; // @[:@133417.4 RegFile.scala 76:16:@133424.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@133423.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@133427.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@133421.4]
  assign regs_397_clock = clock; // @[:@133430.4]
  assign regs_397_reset = io_reset; // @[:@133431.4 RegFile.scala 76:16:@133438.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@133437.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@133441.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@133435.4]
  assign regs_398_clock = clock; // @[:@133444.4]
  assign regs_398_reset = io_reset; // @[:@133445.4 RegFile.scala 76:16:@133452.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@133451.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@133455.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@133449.4]
  assign regs_399_clock = clock; // @[:@133458.4]
  assign regs_399_reset = io_reset; // @[:@133459.4 RegFile.scala 76:16:@133466.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@133465.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@133469.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@133463.4]
  assign regs_400_clock = clock; // @[:@133472.4]
  assign regs_400_reset = io_reset; // @[:@133473.4 RegFile.scala 76:16:@133480.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@133479.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@133483.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@133477.4]
  assign regs_401_clock = clock; // @[:@133486.4]
  assign regs_401_reset = io_reset; // @[:@133487.4 RegFile.scala 76:16:@133494.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@133493.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@133497.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@133491.4]
  assign regs_402_clock = clock; // @[:@133500.4]
  assign regs_402_reset = io_reset; // @[:@133501.4 RegFile.scala 76:16:@133508.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@133507.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@133511.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@133505.4]
  assign regs_403_clock = clock; // @[:@133514.4]
  assign regs_403_reset = io_reset; // @[:@133515.4 RegFile.scala 76:16:@133522.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@133521.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@133525.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@133519.4]
  assign regs_404_clock = clock; // @[:@133528.4]
  assign regs_404_reset = io_reset; // @[:@133529.4 RegFile.scala 76:16:@133536.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@133535.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@133539.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@133533.4]
  assign regs_405_clock = clock; // @[:@133542.4]
  assign regs_405_reset = io_reset; // @[:@133543.4 RegFile.scala 76:16:@133550.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@133549.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@133553.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@133547.4]
  assign regs_406_clock = clock; // @[:@133556.4]
  assign regs_406_reset = io_reset; // @[:@133557.4 RegFile.scala 76:16:@133564.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@133563.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@133567.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@133561.4]
  assign regs_407_clock = clock; // @[:@133570.4]
  assign regs_407_reset = io_reset; // @[:@133571.4 RegFile.scala 76:16:@133578.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@133577.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@133581.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@133575.4]
  assign regs_408_clock = clock; // @[:@133584.4]
  assign regs_408_reset = io_reset; // @[:@133585.4 RegFile.scala 76:16:@133592.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@133591.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@133595.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@133589.4]
  assign regs_409_clock = clock; // @[:@133598.4]
  assign regs_409_reset = io_reset; // @[:@133599.4 RegFile.scala 76:16:@133606.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@133605.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@133609.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@133603.4]
  assign regs_410_clock = clock; // @[:@133612.4]
  assign regs_410_reset = io_reset; // @[:@133613.4 RegFile.scala 76:16:@133620.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@133619.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@133623.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@133617.4]
  assign regs_411_clock = clock; // @[:@133626.4]
  assign regs_411_reset = io_reset; // @[:@133627.4 RegFile.scala 76:16:@133634.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@133633.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@133637.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@133631.4]
  assign regs_412_clock = clock; // @[:@133640.4]
  assign regs_412_reset = io_reset; // @[:@133641.4 RegFile.scala 76:16:@133648.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@133647.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@133651.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@133645.4]
  assign regs_413_clock = clock; // @[:@133654.4]
  assign regs_413_reset = io_reset; // @[:@133655.4 RegFile.scala 76:16:@133662.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@133661.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@133665.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@133659.4]
  assign regs_414_clock = clock; // @[:@133668.4]
  assign regs_414_reset = io_reset; // @[:@133669.4 RegFile.scala 76:16:@133676.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@133675.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@133679.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@133673.4]
  assign regs_415_clock = clock; // @[:@133682.4]
  assign regs_415_reset = io_reset; // @[:@133683.4 RegFile.scala 76:16:@133690.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@133689.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@133693.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@133687.4]
  assign regs_416_clock = clock; // @[:@133696.4]
  assign regs_416_reset = io_reset; // @[:@133697.4 RegFile.scala 76:16:@133704.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@133703.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@133707.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@133701.4]
  assign regs_417_clock = clock; // @[:@133710.4]
  assign regs_417_reset = io_reset; // @[:@133711.4 RegFile.scala 76:16:@133718.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@133717.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@133721.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@133715.4]
  assign regs_418_clock = clock; // @[:@133724.4]
  assign regs_418_reset = io_reset; // @[:@133725.4 RegFile.scala 76:16:@133732.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@133731.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@133735.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@133729.4]
  assign regs_419_clock = clock; // @[:@133738.4]
  assign regs_419_reset = io_reset; // @[:@133739.4 RegFile.scala 76:16:@133746.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@133745.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@133749.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@133743.4]
  assign regs_420_clock = clock; // @[:@133752.4]
  assign regs_420_reset = io_reset; // @[:@133753.4 RegFile.scala 76:16:@133760.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@133759.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@133763.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@133757.4]
  assign regs_421_clock = clock; // @[:@133766.4]
  assign regs_421_reset = io_reset; // @[:@133767.4 RegFile.scala 76:16:@133774.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@133773.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@133777.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@133771.4]
  assign regs_422_clock = clock; // @[:@133780.4]
  assign regs_422_reset = io_reset; // @[:@133781.4 RegFile.scala 76:16:@133788.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@133787.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@133791.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@133785.4]
  assign regs_423_clock = clock; // @[:@133794.4]
  assign regs_423_reset = io_reset; // @[:@133795.4 RegFile.scala 76:16:@133802.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@133801.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@133805.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@133799.4]
  assign regs_424_clock = clock; // @[:@133808.4]
  assign regs_424_reset = io_reset; // @[:@133809.4 RegFile.scala 76:16:@133816.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@133815.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@133819.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@133813.4]
  assign regs_425_clock = clock; // @[:@133822.4]
  assign regs_425_reset = io_reset; // @[:@133823.4 RegFile.scala 76:16:@133830.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@133829.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@133833.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@133827.4]
  assign regs_426_clock = clock; // @[:@133836.4]
  assign regs_426_reset = io_reset; // @[:@133837.4 RegFile.scala 76:16:@133844.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@133843.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@133847.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@133841.4]
  assign regs_427_clock = clock; // @[:@133850.4]
  assign regs_427_reset = io_reset; // @[:@133851.4 RegFile.scala 76:16:@133858.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@133857.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@133861.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@133855.4]
  assign regs_428_clock = clock; // @[:@133864.4]
  assign regs_428_reset = io_reset; // @[:@133865.4 RegFile.scala 76:16:@133872.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@133871.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@133875.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@133869.4]
  assign regs_429_clock = clock; // @[:@133878.4]
  assign regs_429_reset = io_reset; // @[:@133879.4 RegFile.scala 76:16:@133886.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@133885.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@133889.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@133883.4]
  assign regs_430_clock = clock; // @[:@133892.4]
  assign regs_430_reset = io_reset; // @[:@133893.4 RegFile.scala 76:16:@133900.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@133899.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@133903.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@133897.4]
  assign regs_431_clock = clock; // @[:@133906.4]
  assign regs_431_reset = io_reset; // @[:@133907.4 RegFile.scala 76:16:@133914.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@133913.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@133917.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@133911.4]
  assign regs_432_clock = clock; // @[:@133920.4]
  assign regs_432_reset = io_reset; // @[:@133921.4 RegFile.scala 76:16:@133928.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@133927.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@133931.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@133925.4]
  assign regs_433_clock = clock; // @[:@133934.4]
  assign regs_433_reset = io_reset; // @[:@133935.4 RegFile.scala 76:16:@133942.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@133941.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@133945.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@133939.4]
  assign regs_434_clock = clock; // @[:@133948.4]
  assign regs_434_reset = io_reset; // @[:@133949.4 RegFile.scala 76:16:@133956.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@133955.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@133959.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@133953.4]
  assign regs_435_clock = clock; // @[:@133962.4]
  assign regs_435_reset = io_reset; // @[:@133963.4 RegFile.scala 76:16:@133970.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@133969.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@133973.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@133967.4]
  assign regs_436_clock = clock; // @[:@133976.4]
  assign regs_436_reset = io_reset; // @[:@133977.4 RegFile.scala 76:16:@133984.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@133983.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@133987.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@133981.4]
  assign regs_437_clock = clock; // @[:@133990.4]
  assign regs_437_reset = io_reset; // @[:@133991.4 RegFile.scala 76:16:@133998.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@133997.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@134001.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@133995.4]
  assign regs_438_clock = clock; // @[:@134004.4]
  assign regs_438_reset = io_reset; // @[:@134005.4 RegFile.scala 76:16:@134012.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@134011.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@134015.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@134009.4]
  assign regs_439_clock = clock; // @[:@134018.4]
  assign regs_439_reset = io_reset; // @[:@134019.4 RegFile.scala 76:16:@134026.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@134025.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@134029.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@134023.4]
  assign regs_440_clock = clock; // @[:@134032.4]
  assign regs_440_reset = io_reset; // @[:@134033.4 RegFile.scala 76:16:@134040.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@134039.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@134043.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@134037.4]
  assign regs_441_clock = clock; // @[:@134046.4]
  assign regs_441_reset = io_reset; // @[:@134047.4 RegFile.scala 76:16:@134054.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@134053.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@134057.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@134051.4]
  assign regs_442_clock = clock; // @[:@134060.4]
  assign regs_442_reset = io_reset; // @[:@134061.4 RegFile.scala 76:16:@134068.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@134067.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@134071.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@134065.4]
  assign regs_443_clock = clock; // @[:@134074.4]
  assign regs_443_reset = io_reset; // @[:@134075.4 RegFile.scala 76:16:@134082.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@134081.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@134085.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@134079.4]
  assign regs_444_clock = clock; // @[:@134088.4]
  assign regs_444_reset = io_reset; // @[:@134089.4 RegFile.scala 76:16:@134096.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@134095.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@134099.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@134093.4]
  assign regs_445_clock = clock; // @[:@134102.4]
  assign regs_445_reset = io_reset; // @[:@134103.4 RegFile.scala 76:16:@134110.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@134109.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@134113.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@134107.4]
  assign regs_446_clock = clock; // @[:@134116.4]
  assign regs_446_reset = io_reset; // @[:@134117.4 RegFile.scala 76:16:@134124.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@134123.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@134127.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@134121.4]
  assign regs_447_clock = clock; // @[:@134130.4]
  assign regs_447_reset = io_reset; // @[:@134131.4 RegFile.scala 76:16:@134138.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@134137.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@134141.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@134135.4]
  assign regs_448_clock = clock; // @[:@134144.4]
  assign regs_448_reset = io_reset; // @[:@134145.4 RegFile.scala 76:16:@134152.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@134151.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@134155.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@134149.4]
  assign regs_449_clock = clock; // @[:@134158.4]
  assign regs_449_reset = io_reset; // @[:@134159.4 RegFile.scala 76:16:@134166.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@134165.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@134169.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@134163.4]
  assign regs_450_clock = clock; // @[:@134172.4]
  assign regs_450_reset = io_reset; // @[:@134173.4 RegFile.scala 76:16:@134180.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@134179.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@134183.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@134177.4]
  assign regs_451_clock = clock; // @[:@134186.4]
  assign regs_451_reset = io_reset; // @[:@134187.4 RegFile.scala 76:16:@134194.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@134193.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@134197.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@134191.4]
  assign regs_452_clock = clock; // @[:@134200.4]
  assign regs_452_reset = io_reset; // @[:@134201.4 RegFile.scala 76:16:@134208.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@134207.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@134211.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@134205.4]
  assign regs_453_clock = clock; // @[:@134214.4]
  assign regs_453_reset = io_reset; // @[:@134215.4 RegFile.scala 76:16:@134222.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@134221.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@134225.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@134219.4]
  assign regs_454_clock = clock; // @[:@134228.4]
  assign regs_454_reset = io_reset; // @[:@134229.4 RegFile.scala 76:16:@134236.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@134235.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@134239.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@134233.4]
  assign regs_455_clock = clock; // @[:@134242.4]
  assign regs_455_reset = io_reset; // @[:@134243.4 RegFile.scala 76:16:@134250.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@134249.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@134253.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@134247.4]
  assign regs_456_clock = clock; // @[:@134256.4]
  assign regs_456_reset = io_reset; // @[:@134257.4 RegFile.scala 76:16:@134264.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@134263.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@134267.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@134261.4]
  assign regs_457_clock = clock; // @[:@134270.4]
  assign regs_457_reset = io_reset; // @[:@134271.4 RegFile.scala 76:16:@134278.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@134277.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@134281.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@134275.4]
  assign regs_458_clock = clock; // @[:@134284.4]
  assign regs_458_reset = io_reset; // @[:@134285.4 RegFile.scala 76:16:@134292.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@134291.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@134295.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@134289.4]
  assign regs_459_clock = clock; // @[:@134298.4]
  assign regs_459_reset = io_reset; // @[:@134299.4 RegFile.scala 76:16:@134306.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@134305.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@134309.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@134303.4]
  assign regs_460_clock = clock; // @[:@134312.4]
  assign regs_460_reset = io_reset; // @[:@134313.4 RegFile.scala 76:16:@134320.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@134319.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@134323.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@134317.4]
  assign regs_461_clock = clock; // @[:@134326.4]
  assign regs_461_reset = io_reset; // @[:@134327.4 RegFile.scala 76:16:@134334.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@134333.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@134337.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@134331.4]
  assign regs_462_clock = clock; // @[:@134340.4]
  assign regs_462_reset = io_reset; // @[:@134341.4 RegFile.scala 76:16:@134348.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@134347.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@134351.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@134345.4]
  assign regs_463_clock = clock; // @[:@134354.4]
  assign regs_463_reset = io_reset; // @[:@134355.4 RegFile.scala 76:16:@134362.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@134361.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@134365.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@134359.4]
  assign regs_464_clock = clock; // @[:@134368.4]
  assign regs_464_reset = io_reset; // @[:@134369.4 RegFile.scala 76:16:@134376.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@134375.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@134379.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@134373.4]
  assign regs_465_clock = clock; // @[:@134382.4]
  assign regs_465_reset = io_reset; // @[:@134383.4 RegFile.scala 76:16:@134390.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@134389.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@134393.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@134387.4]
  assign regs_466_clock = clock; // @[:@134396.4]
  assign regs_466_reset = io_reset; // @[:@134397.4 RegFile.scala 76:16:@134404.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@134403.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@134407.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@134401.4]
  assign regs_467_clock = clock; // @[:@134410.4]
  assign regs_467_reset = io_reset; // @[:@134411.4 RegFile.scala 76:16:@134418.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@134417.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@134421.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@134415.4]
  assign regs_468_clock = clock; // @[:@134424.4]
  assign regs_468_reset = io_reset; // @[:@134425.4 RegFile.scala 76:16:@134432.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@134431.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@134435.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@134429.4]
  assign regs_469_clock = clock; // @[:@134438.4]
  assign regs_469_reset = io_reset; // @[:@134439.4 RegFile.scala 76:16:@134446.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@134445.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@134449.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@134443.4]
  assign regs_470_clock = clock; // @[:@134452.4]
  assign regs_470_reset = io_reset; // @[:@134453.4 RegFile.scala 76:16:@134460.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@134459.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@134463.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@134457.4]
  assign regs_471_clock = clock; // @[:@134466.4]
  assign regs_471_reset = io_reset; // @[:@134467.4 RegFile.scala 76:16:@134474.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@134473.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@134477.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@134471.4]
  assign regs_472_clock = clock; // @[:@134480.4]
  assign regs_472_reset = io_reset; // @[:@134481.4 RegFile.scala 76:16:@134488.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@134487.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@134491.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@134485.4]
  assign regs_473_clock = clock; // @[:@134494.4]
  assign regs_473_reset = io_reset; // @[:@134495.4 RegFile.scala 76:16:@134502.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@134501.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@134505.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@134499.4]
  assign regs_474_clock = clock; // @[:@134508.4]
  assign regs_474_reset = io_reset; // @[:@134509.4 RegFile.scala 76:16:@134516.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@134515.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@134519.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@134513.4]
  assign regs_475_clock = clock; // @[:@134522.4]
  assign regs_475_reset = io_reset; // @[:@134523.4 RegFile.scala 76:16:@134530.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@134529.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@134533.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@134527.4]
  assign regs_476_clock = clock; // @[:@134536.4]
  assign regs_476_reset = io_reset; // @[:@134537.4 RegFile.scala 76:16:@134544.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@134543.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@134547.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@134541.4]
  assign regs_477_clock = clock; // @[:@134550.4]
  assign regs_477_reset = io_reset; // @[:@134551.4 RegFile.scala 76:16:@134558.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@134557.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@134561.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@134555.4]
  assign regs_478_clock = clock; // @[:@134564.4]
  assign regs_478_reset = io_reset; // @[:@134565.4 RegFile.scala 76:16:@134572.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@134571.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@134575.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@134569.4]
  assign regs_479_clock = clock; // @[:@134578.4]
  assign regs_479_reset = io_reset; // @[:@134579.4 RegFile.scala 76:16:@134586.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@134585.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@134589.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@134583.4]
  assign regs_480_clock = clock; // @[:@134592.4]
  assign regs_480_reset = io_reset; // @[:@134593.4 RegFile.scala 76:16:@134600.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@134599.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@134603.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@134597.4]
  assign regs_481_clock = clock; // @[:@134606.4]
  assign regs_481_reset = io_reset; // @[:@134607.4 RegFile.scala 76:16:@134614.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@134613.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@134617.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@134611.4]
  assign regs_482_clock = clock; // @[:@134620.4]
  assign regs_482_reset = io_reset; // @[:@134621.4 RegFile.scala 76:16:@134628.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@134627.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@134631.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@134625.4]
  assign regs_483_clock = clock; // @[:@134634.4]
  assign regs_483_reset = io_reset; // @[:@134635.4 RegFile.scala 76:16:@134642.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@134641.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@134645.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@134639.4]
  assign regs_484_clock = clock; // @[:@134648.4]
  assign regs_484_reset = io_reset; // @[:@134649.4 RegFile.scala 76:16:@134656.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@134655.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@134659.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@134653.4]
  assign regs_485_clock = clock; // @[:@134662.4]
  assign regs_485_reset = io_reset; // @[:@134663.4 RegFile.scala 76:16:@134670.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@134669.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@134673.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@134667.4]
  assign regs_486_clock = clock; // @[:@134676.4]
  assign regs_486_reset = io_reset; // @[:@134677.4 RegFile.scala 76:16:@134684.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@134683.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@134687.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@134681.4]
  assign regs_487_clock = clock; // @[:@134690.4]
  assign regs_487_reset = io_reset; // @[:@134691.4 RegFile.scala 76:16:@134698.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@134697.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@134701.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@134695.4]
  assign regs_488_clock = clock; // @[:@134704.4]
  assign regs_488_reset = io_reset; // @[:@134705.4 RegFile.scala 76:16:@134712.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@134711.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@134715.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@134709.4]
  assign regs_489_clock = clock; // @[:@134718.4]
  assign regs_489_reset = io_reset; // @[:@134719.4 RegFile.scala 76:16:@134726.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@134725.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@134729.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@134723.4]
  assign regs_490_clock = clock; // @[:@134732.4]
  assign regs_490_reset = io_reset; // @[:@134733.4 RegFile.scala 76:16:@134740.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@134739.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@134743.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@134737.4]
  assign regs_491_clock = clock; // @[:@134746.4]
  assign regs_491_reset = io_reset; // @[:@134747.4 RegFile.scala 76:16:@134754.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@134753.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@134757.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@134751.4]
  assign regs_492_clock = clock; // @[:@134760.4]
  assign regs_492_reset = io_reset; // @[:@134761.4 RegFile.scala 76:16:@134768.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@134767.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@134771.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@134765.4]
  assign regs_493_clock = clock; // @[:@134774.4]
  assign regs_493_reset = io_reset; // @[:@134775.4 RegFile.scala 76:16:@134782.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@134781.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@134785.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@134779.4]
  assign regs_494_clock = clock; // @[:@134788.4]
  assign regs_494_reset = io_reset; // @[:@134789.4 RegFile.scala 76:16:@134796.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@134795.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@134799.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@134793.4]
  assign regs_495_clock = clock; // @[:@134802.4]
  assign regs_495_reset = io_reset; // @[:@134803.4 RegFile.scala 76:16:@134810.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@134809.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@134813.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@134807.4]
  assign regs_496_clock = clock; // @[:@134816.4]
  assign regs_496_reset = io_reset; // @[:@134817.4 RegFile.scala 76:16:@134824.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@134823.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@134827.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@134821.4]
  assign regs_497_clock = clock; // @[:@134830.4]
  assign regs_497_reset = io_reset; // @[:@134831.4 RegFile.scala 76:16:@134838.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@134837.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@134841.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@134835.4]
  assign regs_498_clock = clock; // @[:@134844.4]
  assign regs_498_reset = io_reset; // @[:@134845.4 RegFile.scala 76:16:@134852.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@134851.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@134855.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@134849.4]
  assign regs_499_clock = clock; // @[:@134858.4]
  assign regs_499_reset = io_reset; // @[:@134859.4 RegFile.scala 76:16:@134866.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@134865.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@134869.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@134863.4]
  assign regs_500_clock = clock; // @[:@134872.4]
  assign regs_500_reset = io_reset; // @[:@134873.4 RegFile.scala 76:16:@134880.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@134879.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@134883.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@134877.4]
  assign regs_501_clock = clock; // @[:@134886.4]
  assign regs_501_reset = io_reset; // @[:@134887.4 RegFile.scala 76:16:@134894.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@134893.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@134897.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@134891.4]
  assign regs_502_clock = clock; // @[:@134900.4]
  assign regs_502_reset = io_reset; // @[:@134901.4 RegFile.scala 76:16:@134908.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@134907.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@134911.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@134905.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@135420.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@135421.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@135422.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@135423.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@135424.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@135425.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@135426.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@135427.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@135428.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@135429.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@135430.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@135431.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@135432.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@135433.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@135434.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@135435.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@135436.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@135437.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@135438.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@135439.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@135440.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@135441.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@135442.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@135443.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@135444.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@135445.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@135446.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@135447.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@135448.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@135449.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@135450.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@135451.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@135452.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@135453.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@135454.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@135455.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@135456.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@135457.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@135458.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@135459.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@135460.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@135461.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@135462.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@135463.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@135464.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@135465.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@135466.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@135467.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@135468.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@135469.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@135470.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@135471.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@135472.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@135473.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@135474.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@135475.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@135476.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@135477.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@135478.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@135479.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@135480.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@135481.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@135482.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@135483.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@135484.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@135485.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@135486.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@135487.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@135488.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@135489.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@135490.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@135491.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@135492.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@135493.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@135494.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@135495.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@135496.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@135497.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@135498.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@135499.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@135500.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@135501.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@135502.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@135503.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@135504.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@135505.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@135506.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@135507.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@135508.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@135509.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@135510.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@135511.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@135512.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@135513.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@135514.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@135515.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@135516.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@135517.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@135518.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@135519.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@135520.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@135521.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@135522.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@135523.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@135524.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@135525.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@135526.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@135527.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@135528.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@135529.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@135530.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@135531.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@135532.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@135533.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@135534.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@135535.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@135536.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@135537.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@135538.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@135539.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@135540.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@135541.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@135542.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@135543.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@135544.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@135545.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@135546.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@135547.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@135548.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@135549.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@135550.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@135551.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@135552.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@135553.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@135554.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@135555.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@135556.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@135557.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@135558.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@135559.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@135560.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@135561.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@135562.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@135563.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@135564.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@135565.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@135566.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@135567.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@135568.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@135569.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@135570.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@135571.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@135572.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@135573.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@135574.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@135575.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@135576.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@135577.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@135578.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@135579.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@135580.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@135581.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@135582.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@135583.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@135584.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@135585.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@135586.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@135587.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@135588.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@135589.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@135590.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@135591.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@135592.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@135593.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@135594.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@135595.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@135596.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@135597.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@135598.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@135599.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@135600.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@135601.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@135602.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@135603.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@135604.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@135605.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@135606.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@135607.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@135608.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@135609.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@135610.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@135611.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@135612.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@135613.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@135614.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@135615.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@135616.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@135617.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@135618.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@135619.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@135620.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@135621.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@135622.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@135623.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@135624.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@135625.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@135626.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@135627.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@135628.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@135629.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@135630.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@135631.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@135632.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@135633.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@135634.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@135635.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@135636.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@135637.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@135638.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@135639.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@135640.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@135641.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@135642.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@135643.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@135644.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@135645.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@135646.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@135647.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@135648.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@135649.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@135650.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@135651.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@135652.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@135653.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@135654.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@135655.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@135656.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@135657.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@135658.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@135659.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@135660.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@135661.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@135662.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@135663.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@135664.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@135665.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@135666.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@135667.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@135668.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@135669.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@135670.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@135671.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@135672.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@135673.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@135674.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@135675.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@135676.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@135677.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@135678.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@135679.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@135680.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@135681.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@135682.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@135683.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@135684.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@135685.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@135686.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@135687.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@135688.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@135689.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@135690.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@135691.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@135692.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@135693.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@135694.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@135695.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@135696.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@135697.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@135698.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@135699.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@135700.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@135701.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@135702.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@135703.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@135704.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@135705.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@135706.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@135707.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@135708.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@135709.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@135710.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@135711.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@135712.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@135713.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@135714.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@135715.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@135716.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@135717.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@135718.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@135719.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@135720.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@135721.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@135722.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@135723.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@135724.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@135725.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@135726.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@135727.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@135728.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@135729.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@135730.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@135731.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@135732.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@135733.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@135734.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@135735.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@135736.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@135737.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@135738.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@135739.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@135740.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@135741.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@135742.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@135743.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@135744.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@135745.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@135746.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@135747.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@135748.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@135749.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@135750.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@135751.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@135752.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@135753.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@135754.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@135755.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@135756.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@135757.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@135758.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@135759.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@135760.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@135761.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@135762.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@135763.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@135764.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@135765.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@135766.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@135767.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@135768.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@135769.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@135770.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@135771.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@135772.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@135773.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@135774.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@135775.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@135776.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@135777.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@135778.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@135779.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@135780.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@135781.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@135782.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@135783.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@135784.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@135785.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@135786.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@135787.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@135788.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@135789.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@135790.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@135791.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@135792.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@135793.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@135794.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@135795.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@135796.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@135797.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@135798.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@135799.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@135800.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@135801.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@135802.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@135803.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@135804.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@135805.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@135806.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@135807.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@135808.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@135809.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@135810.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@135811.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@135812.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@135813.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@135814.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@135815.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@135816.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@135817.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@135818.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@135819.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@135820.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@135821.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@135822.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@135823.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@135824.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@135825.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@135826.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@135827.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@135828.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@135829.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@135830.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@135831.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@135832.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@135833.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@135834.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@135835.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@135836.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@135837.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@135838.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@135839.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@135840.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@135841.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@135842.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@135843.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@135844.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@135845.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@135846.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@135847.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@135848.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@135849.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@135850.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@135851.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@135852.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@135853.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@135854.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@135855.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@135856.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@135857.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@135858.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@135859.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@135860.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@135861.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@135862.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@135863.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@135864.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@135865.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@135866.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@135867.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@135868.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@135869.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@135870.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@135871.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@135872.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@135873.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@135874.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@135875.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@135876.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@135877.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@135878.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@135879.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@135880.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@135881.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@135882.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@135883.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@135884.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@135885.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@135886.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@135887.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@135888.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@135889.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@135890.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@135891.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@135892.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@135893.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@135894.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@135895.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@135896.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@135897.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@135898.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@135899.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@135900.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@135901.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@135902.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@135903.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@135904.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@135905.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@135906.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@135907.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@135908.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@135909.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@135910.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@135911.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@135912.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@135913.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@135914.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@135915.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@135916.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@135917.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@135918.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@135919.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@135920.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@135921.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@135922.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@135923.4]
endmodule
module RetimeWrapper_844( // @[:@135947.2]
  input         clock, // @[:@135948.4]
  input         reset, // @[:@135949.4]
  input  [39:0] io_in, // @[:@135950.4]
  output [39:0] io_out // @[:@135950.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@135952.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@135952.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@135952.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@135952.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@135952.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@135952.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@135952.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@135965.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@135964.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@135963.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@135962.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@135961.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@135959.4]
endmodule
module FringeFF_503( // @[:@135967.2]
  input         clock, // @[:@135968.4]
  input         reset, // @[:@135969.4]
  input  [39:0] io_in, // @[:@135970.4]
  output [39:0] io_out, // @[:@135970.4]
  input         io_enable // @[:@135970.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@135973.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@135973.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@135973.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@135973.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@135978.4 package.scala 96:25:@135979.4]
  RetimeWrapper_844 RetimeWrapper ( // @[package.scala 93:22:@135973.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@135978.4 package.scala 96:25:@135979.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@135990.4]
  assign RetimeWrapper_clock = clock; // @[:@135974.4]
  assign RetimeWrapper_reset = reset; // @[:@135975.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@135976.4]
endmodule
module FringeCounter( // @[:@135992.2]
  input   clock, // @[:@135993.4]
  input   reset, // @[:@135994.4]
  input   io_enable, // @[:@135995.4]
  output  io_done // @[:@135995.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@135997.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@135997.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@135997.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@135997.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@135997.4]
  wire [40:0] count; // @[Cat.scala 30:58:@136004.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@136005.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@136006.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@136007.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@136009.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@135997.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@136004.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@136005.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@136006.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@136007.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@136009.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@136020.4]
  assign reg$_clock = clock; // @[:@135998.4]
  assign reg$_reset = reset; // @[:@135999.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@136011.6 FringeCounter.scala 37:15:@136014.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@136002.4]
endmodule
module FringeFF_504( // @[:@136054.2]
  input   clock, // @[:@136055.4]
  input   reset, // @[:@136056.4]
  input   io_in, // @[:@136057.4]
  input   io_reset, // @[:@136057.4]
  output  io_out, // @[:@136057.4]
  input   io_enable // @[:@136057.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@136060.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@136060.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@136060.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@136060.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@136060.4]
  wire  _T_18; // @[package.scala 96:25:@136065.4 package.scala 96:25:@136066.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@136071.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@136060.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@136065.4 package.scala 96:25:@136066.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@136071.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@136077.4]
  assign RetimeWrapper_clock = clock; // @[:@136061.4]
  assign RetimeWrapper_reset = reset; // @[:@136062.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@136064.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@136063.4]
endmodule
module Depulser( // @[:@136079.2]
  input   clock, // @[:@136080.4]
  input   reset, // @[:@136081.4]
  input   io_in, // @[:@136082.4]
  input   io_rst, // @[:@136082.4]
  output  io_out // @[:@136082.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@136084.4]
  wire  r_reset; // @[Depulser.scala 14:17:@136084.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@136084.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@136084.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@136084.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@136084.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@136084.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@136093.4]
  assign r_clock = clock; // @[:@136085.4]
  assign r_reset = reset; // @[:@136086.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@136088.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@136092.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@136091.4]
endmodule
module Fringe( // @[:@136095.2]
  input         clock, // @[:@136096.4]
  input         reset, // @[:@136097.4]
  input  [31:0] io_raddr, // @[:@136098.4]
  input         io_wen, // @[:@136098.4]
  input  [31:0] io_waddr, // @[:@136098.4]
  input  [63:0] io_wdata, // @[:@136098.4]
  output [63:0] io_rdata, // @[:@136098.4]
  output        io_enable, // @[:@136098.4]
  input         io_done, // @[:@136098.4]
  output        io_reset, // @[:@136098.4]
  output [63:0] io_argIns_0, // @[:@136098.4]
  output [63:0] io_argIns_1, // @[:@136098.4]
  input         io_argOuts_0_valid, // @[:@136098.4]
  input  [63:0] io_argOuts_0_bits, // @[:@136098.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@136098.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@136098.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@136098.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@136098.4]
  output        io_memStreams_stores_0_data_ready, // @[:@136098.4]
  input         io_memStreams_stores_0_data_valid, // @[:@136098.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@136098.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@136098.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@136098.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@136098.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@136098.4]
  input         io_dram_0_cmd_ready, // @[:@136098.4]
  output        io_dram_0_cmd_valid, // @[:@136098.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@136098.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@136098.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@136098.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@136098.4]
  input         io_dram_0_wdata_ready, // @[:@136098.4]
  output        io_dram_0_wdata_valid, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@136098.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@136098.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@136098.4]
  output        io_dram_0_rresp_ready, // @[:@136098.4]
  output        io_dram_0_wresp_ready, // @[:@136098.4]
  input         io_dram_0_wresp_valid, // @[:@136098.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@136098.4]
  input         io_dram_1_cmd_ready, // @[:@136098.4]
  output        io_dram_1_cmd_valid, // @[:@136098.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@136098.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@136098.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@136098.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@136098.4]
  input         io_dram_1_wdata_ready, // @[:@136098.4]
  output        io_dram_1_wdata_valid, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@136098.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@136098.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@136098.4]
  output        io_dram_1_rresp_ready, // @[:@136098.4]
  output        io_dram_1_wresp_ready, // @[:@136098.4]
  input         io_dram_1_wresp_valid, // @[:@136098.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@136098.4]
  input         io_dram_2_cmd_ready, // @[:@136098.4]
  output        io_dram_2_cmd_valid, // @[:@136098.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@136098.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@136098.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@136098.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@136098.4]
  input         io_dram_2_wdata_ready, // @[:@136098.4]
  output        io_dram_2_wdata_valid, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@136098.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@136098.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@136098.4]
  output        io_dram_2_rresp_ready, // @[:@136098.4]
  output        io_dram_2_wresp_ready, // @[:@136098.4]
  input         io_dram_2_wresp_valid, // @[:@136098.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@136098.4]
  input         io_dram_3_cmd_ready, // @[:@136098.4]
  output        io_dram_3_cmd_valid, // @[:@136098.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@136098.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@136098.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@136098.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@136098.4]
  input         io_dram_3_wdata_ready, // @[:@136098.4]
  output        io_dram_3_wdata_valid, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@136098.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@136098.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@136098.4]
  output        io_dram_3_rresp_ready, // @[:@136098.4]
  output        io_dram_3_wresp_ready, // @[:@136098.4]
  input         io_dram_3_wresp_valid, // @[:@136098.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@136098.4]
  input         io_heap_0_req_valid, // @[:@136098.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@136098.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@136098.4]
  output        io_heap_0_resp_valid, // @[:@136098.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@136098.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@136098.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@136104.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@136104.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@136104.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@136104.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@137097.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@137097.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@137097.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@138057.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@138057.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@138057.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@139017.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@139017.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@139017.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@139017.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@139977.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@139977.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@139977.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@139977.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@139977.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@139977.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@139977.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@139977.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@139977.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@139977.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@139977.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@139977.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@139986.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@139986.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@139986.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@139986.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@139986.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@139986.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@139986.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@139986.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@139986.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@142036.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@142036.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@142036.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@142036.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@142055.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@142055.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@142055.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@142055.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@142055.4]
  wire [63:0] _T_1020; // @[:@142013.4 :@142014.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@142015.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@142017.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@142019.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@142021.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@142023.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@142025.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@142027.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@142063.4]
  reg  _T_1047; // @[package.scala 152:20:@142066.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@142068.4]
  wire  _T_1049; // @[package.scala 153:8:@142069.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@142073.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@142074.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@142077.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@142078.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@142080.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@142081.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@142083.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@142086.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@142065.4 Fringe.scala 163:24:@142084.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@142065.4 Fringe.scala 162:28:@142082.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@142087.4]
  wire  alloc; // @[Fringe.scala 202:38:@143717.4]
  wire  dealloc; // @[Fringe.scala 203:40:@143718.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@143719.4]
  reg  _T_1572; // @[package.scala 152:20:@143720.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@143722.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@136104.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@137097.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@138057.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@139017.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@139977.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@139986.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@142036.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@142055.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@142013.4 :@142014.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@142015.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@142017.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@142019.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@142021.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@142023.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@142025.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@142027.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@142063.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@142068.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@142069.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@142073.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@142074.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@142077.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@142078.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@142080.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@142081.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@142083.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@142086.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@142065.4 Fringe.scala 163:24:@142084.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@142065.4 Fringe.scala 162:28:@142082.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@142087.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@143717.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@143718.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@143719.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@143722.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@142011.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@142031.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@142032.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@142053.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@142054.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@137023.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@137019.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@137014.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@137013.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@143215.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@143214.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@143213.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@143211.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@143210.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@143208.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@143192.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@143193.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@143194.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@143195.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@143196.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@143197.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@143198.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@143199.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@143200.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@143201.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@143202.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@143203.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@143204.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@143205.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@143206.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@143207.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@143128.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@143129.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@143130.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@143131.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@143132.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@143133.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@143134.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@143135.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@143136.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@143137.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@143138.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@143139.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@143140.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@143141.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@143142.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@143143.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@143144.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@143145.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@143146.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@143147.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@143148.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@143149.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@143150.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@143151.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@143152.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@143153.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@143154.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@143155.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@143156.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@143157.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@143158.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@143159.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@143160.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@143161.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@143162.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@143163.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@143164.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@143165.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@143166.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@143167.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@143168.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@143169.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@143170.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@143171.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@143172.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@143173.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@143174.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@143175.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@143176.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@143177.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@143178.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@143179.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@143180.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@143181.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@143182.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@143183.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@143184.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@143185.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@143186.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@143187.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@143188.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@143189.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@143190.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@143191.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@143127.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@143126.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@143107.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@143327.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@143326.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@143325.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@143323.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@143322.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@143320.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@143304.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@143305.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@143306.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@143307.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@143308.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@143309.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@143310.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@143311.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@143312.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@143313.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@143314.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@143315.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@143316.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@143317.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@143318.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@143319.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@143240.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@143241.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@143242.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@143243.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@143244.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@143245.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@143246.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@143247.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@143248.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@143249.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@143250.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@143251.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@143252.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@143253.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@143254.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@143255.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@143256.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@143257.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@143258.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@143259.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@143260.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@143261.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@143262.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@143263.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@143264.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@143265.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@143266.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@143267.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@143268.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@143269.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@143270.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@143271.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@143272.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@143273.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@143274.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@143275.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@143276.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@143277.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@143278.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@143279.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@143280.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@143281.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@143282.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@143283.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@143284.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@143285.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@143286.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@143287.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@143288.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@143289.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@143290.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@143291.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@143292.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@143293.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@143294.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@143295.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@143296.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@143297.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@143298.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@143299.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@143300.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@143301.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@143302.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@143303.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@143239.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@143238.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@143219.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@143439.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@143438.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@143437.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@143435.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@143434.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@143432.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@143416.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@143417.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@143418.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@143419.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@143420.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@143421.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@143422.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@143423.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@143424.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@143425.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@143426.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@143427.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@143428.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@143429.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@143430.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@143431.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@143352.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@143353.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@143354.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@143355.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@143356.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@143357.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@143358.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@143359.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@143360.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@143361.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@143362.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@143363.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@143364.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@143365.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@143366.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@143367.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@143368.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@143369.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@143370.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@143371.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@143372.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@143373.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@143374.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@143375.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@143376.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@143377.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@143378.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@143379.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@143380.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@143381.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@143382.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@143383.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@143384.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@143385.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@143386.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@143387.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@143388.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@143389.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@143390.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@143391.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@143392.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@143393.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@143394.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@143395.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@143396.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@143397.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@143398.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@143399.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@143400.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@143401.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@143402.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@143403.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@143404.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@143405.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@143406.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@143407.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@143408.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@143409.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@143410.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@143411.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@143412.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@143413.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@143414.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@143415.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@143351.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@143350.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@143331.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@143551.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@143550.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@143549.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@143547.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@143546.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@143544.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@143528.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@143529.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@143530.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@143531.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@143532.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@143533.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@143534.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@143535.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@143536.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@143537.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@143538.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@143539.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@143540.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@143541.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@143542.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@143543.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@143464.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@143465.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@143466.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@143467.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@143468.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@143469.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@143470.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@143471.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@143472.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@143473.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@143474.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@143475.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@143476.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@143477.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@143478.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@143479.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@143480.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@143481.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@143482.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@143483.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@143484.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@143485.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@143486.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@143487.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@143488.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@143489.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@143490.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@143491.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@143492.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@143493.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@143494.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@143495.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@143496.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@143497.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@143498.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@143499.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@143500.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@143501.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@143502.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@143503.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@143504.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@143505.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@143506.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@143507.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@143508.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@143509.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@143510.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@143511.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@143512.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@143513.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@143514.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@143515.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@143516.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@143517.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@143518.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@143519.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@143520.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@143521.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@143522.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@143523.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@143524.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@143525.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@143526.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@143527.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@143463.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@143462.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@143443.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@139982.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@139981.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@139980.4]
  assign dramArbs_0_clock = clock; // @[:@136105.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@136106.4 Fringe.scala 187:30:@143097.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@143101.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@137022.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@137021.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@137020.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@137018.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@137017.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@137016.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@137015.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@143216.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@143209.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@143106.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@143105.4]
  assign dramArbs_1_clock = clock; // @[:@137098.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@137099.4 Fringe.scala 187:30:@143098.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@143102.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@143328.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@143321.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@143218.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@143217.4]
  assign dramArbs_2_clock = clock; // @[:@138058.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@138059.4 Fringe.scala 187:30:@143099.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@143103.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@143440.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@143433.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@143330.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@143329.4]
  assign dramArbs_3_clock = clock; // @[:@139018.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@139019.4 Fringe.scala 187:30:@143100.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@143104.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@143552.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@143545.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@143442.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@143441.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@139985.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@139984.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@139983.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@143724.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@143725.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@143726.4]
  assign regs_clock = clock; // @[:@139987.4]
  assign regs_reset = reset; // @[:@139988.4 Fringe.scala 139:14:@142035.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@142007.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@142009.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@142008.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@142010.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@142033.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@142085.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@142089.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@142092.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@142091.4]
  assign timeoutCtr_clock = clock; // @[:@142037.4]
  assign timeoutCtr_reset = reset; // @[:@142038.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@142052.4]
  assign depulser_clock = clock; // @[:@142056.4]
  assign depulser_reset = reset; // @[:@142057.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@142062.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@142064.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@143741.2]
  input         clock, // @[:@143742.4]
  input         reset, // @[:@143743.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@143744.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@143744.4]
  input         io_S_AXI_AWVALID, // @[:@143744.4]
  output        io_S_AXI_AWREADY, // @[:@143744.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@143744.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@143744.4]
  input         io_S_AXI_ARVALID, // @[:@143744.4]
  output        io_S_AXI_ARREADY, // @[:@143744.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@143744.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@143744.4]
  input         io_S_AXI_WVALID, // @[:@143744.4]
  output        io_S_AXI_WREADY, // @[:@143744.4]
  output [31:0] io_S_AXI_RDATA, // @[:@143744.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@143744.4]
  output        io_S_AXI_RVALID, // @[:@143744.4]
  input         io_S_AXI_RREADY, // @[:@143744.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@143744.4]
  output        io_S_AXI_BVALID, // @[:@143744.4]
  input         io_S_AXI_BREADY, // @[:@143744.4]
  output [31:0] io_raddr, // @[:@143744.4]
  output        io_wen, // @[:@143744.4]
  output [31:0] io_waddr, // @[:@143744.4]
  output [31:0] io_wdata, // @[:@143744.4]
  input  [31:0] io_rdata // @[:@143744.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@143746.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@143770.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@143766.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@143762.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@143761.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@143760.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@143759.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@143757.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@143756.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@143778.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@143781.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@143779.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@143780.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@143782.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@143777.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@143774.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@143773.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@143772.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@143771.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@143769.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@143768.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@143767.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@143765.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@143764.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@143763.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@143758.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@143755.4]
endmodule
module MAGToAXI4Bridge( // @[:@143784.2]
  output         io_in_cmd_ready, // @[:@143787.4]
  input          io_in_cmd_valid, // @[:@143787.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@143787.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@143787.4]
  input          io_in_cmd_bits_isWr, // @[:@143787.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@143787.4]
  output         io_in_wdata_ready, // @[:@143787.4]
  input          io_in_wdata_valid, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@143787.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@143787.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@143787.4]
  input          io_in_wdata_bits_wlast, // @[:@143787.4]
  input          io_in_rresp_ready, // @[:@143787.4]
  input          io_in_wresp_ready, // @[:@143787.4]
  output         io_in_wresp_valid, // @[:@143787.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@143787.4]
  output [31:0]  io_M_AXI_AWID, // @[:@143787.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@143787.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@143787.4]
  output         io_M_AXI_AWVALID, // @[:@143787.4]
  input          io_M_AXI_AWREADY, // @[:@143787.4]
  output [31:0]  io_M_AXI_ARID, // @[:@143787.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@143787.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@143787.4]
  output         io_M_AXI_ARVALID, // @[:@143787.4]
  input          io_M_AXI_ARREADY, // @[:@143787.4]
  output [511:0] io_M_AXI_WDATA, // @[:@143787.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@143787.4]
  output         io_M_AXI_WLAST, // @[:@143787.4]
  output         io_M_AXI_WVALID, // @[:@143787.4]
  input          io_M_AXI_WREADY, // @[:@143787.4]
  output         io_M_AXI_RREADY, // @[:@143787.4]
  input  [31:0]  io_M_AXI_BID, // @[:@143787.4]
  input          io_M_AXI_BVALID, // @[:@143787.4]
  output         io_M_AXI_BREADY // @[:@143787.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@143944.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@143945.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@143946.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@143954.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@143981.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@143986.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@143997.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@144006.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@144015.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@144024.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@144033.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@144042.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@144050.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@143944.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@143945.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@143946.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@143954.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@143981.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@143986.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@143997.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@144006.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@144015.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@144024.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@144033.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@144042.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@144050.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@143958.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@144055.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@144108.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@144110.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@143959.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@143960.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@143964.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@143972.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@143942.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@143943.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@143947.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@143956.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@143988.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@144052.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@144053.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@144054.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@144105.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@144106.4]
endmodule
module FringeZynq( // @[:@145096.2]
  input          clock, // @[:@145097.4]
  input          reset, // @[:@145098.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@145099.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@145099.4]
  input          io_S_AXI_AWVALID, // @[:@145099.4]
  output         io_S_AXI_AWREADY, // @[:@145099.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@145099.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@145099.4]
  input          io_S_AXI_ARVALID, // @[:@145099.4]
  output         io_S_AXI_ARREADY, // @[:@145099.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@145099.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@145099.4]
  input          io_S_AXI_WVALID, // @[:@145099.4]
  output         io_S_AXI_WREADY, // @[:@145099.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@145099.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@145099.4]
  output         io_S_AXI_RVALID, // @[:@145099.4]
  input          io_S_AXI_RREADY, // @[:@145099.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@145099.4]
  output         io_S_AXI_BVALID, // @[:@145099.4]
  input          io_S_AXI_BREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@145099.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@145099.4]
  output         io_M_AXI_0_AWVALID, // @[:@145099.4]
  input          io_M_AXI_0_AWREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@145099.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@145099.4]
  output         io_M_AXI_0_ARVALID, // @[:@145099.4]
  input          io_M_AXI_0_ARREADY, // @[:@145099.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@145099.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@145099.4]
  output         io_M_AXI_0_WLAST, // @[:@145099.4]
  output         io_M_AXI_0_WVALID, // @[:@145099.4]
  input          io_M_AXI_0_WREADY, // @[:@145099.4]
  output         io_M_AXI_0_RREADY, // @[:@145099.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@145099.4]
  input          io_M_AXI_0_BVALID, // @[:@145099.4]
  output         io_M_AXI_0_BREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@145099.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@145099.4]
  output         io_M_AXI_1_AWVALID, // @[:@145099.4]
  input          io_M_AXI_1_AWREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@145099.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@145099.4]
  output         io_M_AXI_1_ARVALID, // @[:@145099.4]
  input          io_M_AXI_1_ARREADY, // @[:@145099.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@145099.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@145099.4]
  output         io_M_AXI_1_WLAST, // @[:@145099.4]
  output         io_M_AXI_1_WVALID, // @[:@145099.4]
  input          io_M_AXI_1_WREADY, // @[:@145099.4]
  output         io_M_AXI_1_RREADY, // @[:@145099.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@145099.4]
  input          io_M_AXI_1_BVALID, // @[:@145099.4]
  output         io_M_AXI_1_BREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@145099.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@145099.4]
  output         io_M_AXI_2_AWVALID, // @[:@145099.4]
  input          io_M_AXI_2_AWREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@145099.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@145099.4]
  output         io_M_AXI_2_ARVALID, // @[:@145099.4]
  input          io_M_AXI_2_ARREADY, // @[:@145099.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@145099.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@145099.4]
  output         io_M_AXI_2_WLAST, // @[:@145099.4]
  output         io_M_AXI_2_WVALID, // @[:@145099.4]
  input          io_M_AXI_2_WREADY, // @[:@145099.4]
  output         io_M_AXI_2_RREADY, // @[:@145099.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@145099.4]
  input          io_M_AXI_2_BVALID, // @[:@145099.4]
  output         io_M_AXI_2_BREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@145099.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@145099.4]
  output         io_M_AXI_3_AWVALID, // @[:@145099.4]
  input          io_M_AXI_3_AWREADY, // @[:@145099.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@145099.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@145099.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@145099.4]
  output         io_M_AXI_3_ARVALID, // @[:@145099.4]
  input          io_M_AXI_3_ARREADY, // @[:@145099.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@145099.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@145099.4]
  output         io_M_AXI_3_WLAST, // @[:@145099.4]
  output         io_M_AXI_3_WVALID, // @[:@145099.4]
  input          io_M_AXI_3_WREADY, // @[:@145099.4]
  output         io_M_AXI_3_RREADY, // @[:@145099.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@145099.4]
  input          io_M_AXI_3_BVALID, // @[:@145099.4]
  output         io_M_AXI_3_BREADY, // @[:@145099.4]
  output         io_enable, // @[:@145099.4]
  input          io_done, // @[:@145099.4]
  output         io_reset, // @[:@145099.4]
  output [63:0]  io_argIns_0, // @[:@145099.4]
  output [63:0]  io_argIns_1, // @[:@145099.4]
  input          io_argOuts_0_valid, // @[:@145099.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@145099.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@145099.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@145099.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@145099.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@145099.4]
  output         io_memStreams_stores_0_data_ready, // @[:@145099.4]
  input          io_memStreams_stores_0_data_valid, // @[:@145099.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@145099.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@145099.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@145099.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@145099.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@145099.4]
  input          io_heap_0_req_valid, // @[:@145099.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@145099.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@145099.4]
  output         io_heap_0_resp_valid, // @[:@145099.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@145099.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@145099.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@145570.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@145570.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@145570.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@146476.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@146476.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@146476.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@146476.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@146476.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@146476.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@146476.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@146476.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@146626.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@146626.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@146626.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@146626.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@146626.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@146626.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@146626.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@146782.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@146782.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@146782.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@146782.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@146782.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@146782.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@146782.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@146938.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@146938.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@146938.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@146938.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@146938.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@146938.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@146938.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@147094.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@147094.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@147094.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@147094.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@147094.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@147094.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@147094.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@147094.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@145570.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@146476.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@146626.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@146782.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@146938.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@147094.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@146494.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@146490.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@146486.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@146485.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@146484.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@146483.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@146481.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@146480.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@146781.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@146779.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@146778.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@146771.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@146769.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@146767.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@146766.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@146759.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@146757.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@146756.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@146755.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@146754.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@146746.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@146741.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@146937.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@146935.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@146934.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@146927.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@146925.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@146923.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@146922.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@146915.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@146913.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@146912.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@146911.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@146910.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@146902.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@146897.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@147093.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@147091.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@147090.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@147083.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@147081.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@147079.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@147078.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@147071.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@147069.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@147068.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@147067.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@147066.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@147058.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@147053.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@147249.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@147247.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@147246.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@147239.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@147237.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@147235.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@147234.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@147227.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@147225.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@147224.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@147223.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@147222.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@147214.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@147209.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@146504.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@146508.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@146509.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@146510.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@146597.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@146593.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@146588.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@146587.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@146622.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@146621.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@146620.4]
  assign fringeCommon_clock = clock; // @[:@145571.4]
  assign fringeCommon_reset = reset; // @[:@145572.4 FringeZynq.scala 117:22:@146507.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@146498.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@146499.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@146500.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@146501.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@146505.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@146512.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@146511.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@146596.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@146595.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@146594.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@146592.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@146591.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@146590.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@146589.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@146740.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@146733.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@146630.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@146629.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@146896.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@146889.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@146786.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@146785.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@147052.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@147045.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@146942.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@146941.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@147208.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@147201.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@147098.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@147097.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@146625.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@146624.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@146623.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@146477.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@146478.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@146497.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@146496.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@146495.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@146493.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@146492.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@146491.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@146489.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@146488.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@146487.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@146482.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@146479.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@146502.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@146739.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@146738.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@146737.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@146735.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@146734.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@146732.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@146716.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@146717.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@146718.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@146719.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@146720.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@146721.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@146722.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@146723.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@146724.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@146725.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@146726.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@146727.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@146728.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@146729.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@146730.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@146731.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@146652.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@146653.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@146654.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@146655.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@146656.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@146657.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@146658.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@146659.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@146660.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@146661.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@146662.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@146663.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@146664.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@146665.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@146666.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@146667.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@146668.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@146669.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@146670.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@146671.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@146672.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@146673.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@146674.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@146675.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@146676.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@146677.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@146678.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@146679.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@146680.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@146681.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@146682.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@146683.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@146684.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@146685.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@146686.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@146687.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@146688.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@146689.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@146690.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@146691.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@146692.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@146693.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@146694.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@146695.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@146696.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@146697.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@146698.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@146699.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@146700.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@146701.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@146702.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@146703.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@146704.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@146705.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@146706.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@146707.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@146708.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@146709.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@146710.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@146711.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@146712.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@146713.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@146714.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@146715.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@146651.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@146650.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@146631.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@146770.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@146758.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@146753.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@146745.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@146742.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@146895.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@146894.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@146893.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@146891.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@146890.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@146888.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@146872.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@146873.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@146874.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@146875.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@146876.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@146877.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@146878.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@146879.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@146880.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@146881.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@146882.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@146883.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@146884.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@146885.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@146886.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@146887.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@146808.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@146809.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@146810.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@146811.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@146812.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@146813.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@146814.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@146815.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@146816.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@146817.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@146818.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@146819.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@146820.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@146821.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@146822.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@146823.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@146824.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@146825.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@146826.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@146827.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@146828.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@146829.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@146830.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@146831.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@146832.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@146833.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@146834.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@146835.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@146836.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@146837.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@146838.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@146839.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@146840.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@146841.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@146842.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@146843.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@146844.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@146845.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@146846.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@146847.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@146848.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@146849.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@146850.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@146851.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@146852.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@146853.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@146854.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@146855.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@146856.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@146857.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@146858.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@146859.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@146860.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@146861.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@146862.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@146863.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@146864.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@146865.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@146866.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@146867.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@146868.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@146869.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@146870.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@146871.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@146807.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@146806.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@146787.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@146926.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@146914.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@146909.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@146901.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@146898.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@147051.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@147050.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@147049.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@147047.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@147046.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@147044.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@147028.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@147029.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@147030.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@147031.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@147032.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@147033.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@147034.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@147035.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@147036.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@147037.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@147038.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@147039.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@147040.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@147041.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@147042.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@147043.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@146964.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@146965.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@146966.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@146967.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@146968.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@146969.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@146970.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@146971.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@146972.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@146973.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@146974.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@146975.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@146976.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@146977.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@146978.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@146979.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@146980.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@146981.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@146982.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@146983.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@146984.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@146985.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@146986.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@146987.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@146988.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@146989.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@146990.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@146991.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@146992.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@146993.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@146994.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@146995.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@146996.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@146997.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@146998.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@146999.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@147000.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@147001.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@147002.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@147003.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@147004.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@147005.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@147006.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@147007.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@147008.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@147009.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@147010.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@147011.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@147012.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@147013.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@147014.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@147015.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@147016.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@147017.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@147018.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@147019.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@147020.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@147021.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@147022.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@147023.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@147024.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@147025.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@147026.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@147027.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@146963.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@146962.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@146943.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@147082.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@147070.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@147065.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@147057.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@147054.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@147207.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@147206.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@147205.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@147203.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@147202.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@147200.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@147184.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@147185.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@147186.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@147187.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@147188.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@147189.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@147190.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@147191.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@147192.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@147193.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@147194.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@147195.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@147196.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@147197.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@147198.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@147199.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@147120.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@147121.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@147122.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@147123.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@147124.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@147125.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@147126.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@147127.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@147128.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@147129.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@147130.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@147131.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@147132.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@147133.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@147134.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@147135.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@147136.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@147137.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@147138.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@147139.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@147140.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@147141.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@147142.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@147143.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@147144.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@147145.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@147146.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@147147.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@147148.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@147149.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@147150.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@147151.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@147152.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@147153.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@147154.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@147155.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@147156.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@147157.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@147158.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@147159.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@147160.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@147161.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@147162.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@147163.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@147164.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@147165.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@147166.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@147167.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@147168.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@147169.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@147170.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@147171.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@147172.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@147173.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@147174.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@147175.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@147176.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@147177.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@147178.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@147179.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@147180.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@147181.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@147182.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@147183.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@147119.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@147118.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@147099.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@147238.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@147226.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@147221.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@147213.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@147210.4]
endmodule
module SpatialIP( // @[:@147251.2]
  input          clock, // @[:@147252.4]
  input          reset, // @[:@147253.4]
  input          io_raddr, // @[:@147254.4]
  input          io_wen, // @[:@147254.4]
  input          io_waddr, // @[:@147254.4]
  input          io_wdata, // @[:@147254.4]
  output         io_rdata, // @[:@147254.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@147254.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@147254.4]
  input          io_S_AXI_AWVALID, // @[:@147254.4]
  output         io_S_AXI_AWREADY, // @[:@147254.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@147254.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@147254.4]
  input          io_S_AXI_ARVALID, // @[:@147254.4]
  output         io_S_AXI_ARREADY, // @[:@147254.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@147254.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@147254.4]
  input          io_S_AXI_WVALID, // @[:@147254.4]
  output         io_S_AXI_WREADY, // @[:@147254.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@147254.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@147254.4]
  output         io_S_AXI_RVALID, // @[:@147254.4]
  input          io_S_AXI_RREADY, // @[:@147254.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@147254.4]
  output         io_S_AXI_BVALID, // @[:@147254.4]
  input          io_S_AXI_BREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@147254.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@147254.4]
  output         io_M_AXI_0_AWLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@147254.4]
  output         io_M_AXI_0_AWVALID, // @[:@147254.4]
  input          io_M_AXI_0_AWREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@147254.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@147254.4]
  output         io_M_AXI_0_ARLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@147254.4]
  output         io_M_AXI_0_ARVALID, // @[:@147254.4]
  input          io_M_AXI_0_ARREADY, // @[:@147254.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@147254.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@147254.4]
  output         io_M_AXI_0_WLAST, // @[:@147254.4]
  output         io_M_AXI_0_WVALID, // @[:@147254.4]
  input          io_M_AXI_0_WREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@147254.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@147254.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@147254.4]
  input          io_M_AXI_0_RLAST, // @[:@147254.4]
  input          io_M_AXI_0_RVALID, // @[:@147254.4]
  output         io_M_AXI_0_RREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@147254.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@147254.4]
  input          io_M_AXI_0_BVALID, // @[:@147254.4]
  output         io_M_AXI_0_BREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@147254.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@147254.4]
  output         io_M_AXI_1_AWLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@147254.4]
  output         io_M_AXI_1_AWVALID, // @[:@147254.4]
  input          io_M_AXI_1_AWREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@147254.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@147254.4]
  output         io_M_AXI_1_ARLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@147254.4]
  output         io_M_AXI_1_ARVALID, // @[:@147254.4]
  input          io_M_AXI_1_ARREADY, // @[:@147254.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@147254.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@147254.4]
  output         io_M_AXI_1_WLAST, // @[:@147254.4]
  output         io_M_AXI_1_WVALID, // @[:@147254.4]
  input          io_M_AXI_1_WREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@147254.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@147254.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@147254.4]
  input          io_M_AXI_1_RLAST, // @[:@147254.4]
  input          io_M_AXI_1_RVALID, // @[:@147254.4]
  output         io_M_AXI_1_RREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@147254.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@147254.4]
  input          io_M_AXI_1_BVALID, // @[:@147254.4]
  output         io_M_AXI_1_BREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@147254.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@147254.4]
  output         io_M_AXI_2_AWLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@147254.4]
  output         io_M_AXI_2_AWVALID, // @[:@147254.4]
  input          io_M_AXI_2_AWREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@147254.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@147254.4]
  output         io_M_AXI_2_ARLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@147254.4]
  output         io_M_AXI_2_ARVALID, // @[:@147254.4]
  input          io_M_AXI_2_ARREADY, // @[:@147254.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@147254.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@147254.4]
  output         io_M_AXI_2_WLAST, // @[:@147254.4]
  output         io_M_AXI_2_WVALID, // @[:@147254.4]
  input          io_M_AXI_2_WREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@147254.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@147254.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@147254.4]
  input          io_M_AXI_2_RLAST, // @[:@147254.4]
  input          io_M_AXI_2_RVALID, // @[:@147254.4]
  output         io_M_AXI_2_RREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@147254.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@147254.4]
  input          io_M_AXI_2_BVALID, // @[:@147254.4]
  output         io_M_AXI_2_BREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@147254.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@147254.4]
  output         io_M_AXI_3_AWLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@147254.4]
  output         io_M_AXI_3_AWVALID, // @[:@147254.4]
  input          io_M_AXI_3_AWREADY, // @[:@147254.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@147254.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@147254.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@147254.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@147254.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@147254.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@147254.4]
  output         io_M_AXI_3_ARLOCK, // @[:@147254.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@147254.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@147254.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@147254.4]
  output         io_M_AXI_3_ARVALID, // @[:@147254.4]
  input          io_M_AXI_3_ARREADY, // @[:@147254.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@147254.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@147254.4]
  output         io_M_AXI_3_WLAST, // @[:@147254.4]
  output         io_M_AXI_3_WVALID, // @[:@147254.4]
  input          io_M_AXI_3_WREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@147254.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@147254.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@147254.4]
  input          io_M_AXI_3_RLAST, // @[:@147254.4]
  input          io_M_AXI_3_RVALID, // @[:@147254.4]
  output         io_M_AXI_3_RREADY, // @[:@147254.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@147254.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@147254.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@147254.4]
  input          io_M_AXI_3_BVALID, // @[:@147254.4]
  output         io_M_AXI_3_BREADY, // @[:@147254.4]
  input          io_TOP_AXI_AWID, // @[:@147254.4]
  input          io_TOP_AXI_AWUSER, // @[:@147254.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@147254.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@147254.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@147254.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@147254.4]
  input          io_TOP_AXI_AWLOCK, // @[:@147254.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@147254.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@147254.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@147254.4]
  input          io_TOP_AXI_AWVALID, // @[:@147254.4]
  input          io_TOP_AXI_AWREADY, // @[:@147254.4]
  input          io_TOP_AXI_ARID, // @[:@147254.4]
  input          io_TOP_AXI_ARUSER, // @[:@147254.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@147254.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@147254.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@147254.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@147254.4]
  input          io_TOP_AXI_ARLOCK, // @[:@147254.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@147254.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@147254.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@147254.4]
  input          io_TOP_AXI_ARVALID, // @[:@147254.4]
  input          io_TOP_AXI_ARREADY, // @[:@147254.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@147254.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@147254.4]
  input          io_TOP_AXI_WLAST, // @[:@147254.4]
  input          io_TOP_AXI_WVALID, // @[:@147254.4]
  input          io_TOP_AXI_WREADY, // @[:@147254.4]
  input          io_TOP_AXI_RID, // @[:@147254.4]
  input          io_TOP_AXI_RUSER, // @[:@147254.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@147254.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@147254.4]
  input          io_TOP_AXI_RLAST, // @[:@147254.4]
  input          io_TOP_AXI_RVALID, // @[:@147254.4]
  input          io_TOP_AXI_RREADY, // @[:@147254.4]
  input          io_TOP_AXI_BID, // @[:@147254.4]
  input          io_TOP_AXI_BUSER, // @[:@147254.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@147254.4]
  input          io_TOP_AXI_BVALID, // @[:@147254.4]
  input          io_TOP_AXI_BREADY, // @[:@147254.4]
  input          io_DWIDTH_AXI_AWID, // @[:@147254.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@147254.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@147254.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@147254.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@147254.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@147254.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@147254.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@147254.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@147254.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@147254.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@147254.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@147254.4]
  input          io_DWIDTH_AXI_ARID, // @[:@147254.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@147254.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@147254.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@147254.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@147254.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@147254.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@147254.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@147254.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@147254.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@147254.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@147254.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@147254.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@147254.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@147254.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@147254.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@147254.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@147254.4]
  input          io_DWIDTH_AXI_RID, // @[:@147254.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@147254.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@147254.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@147254.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@147254.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@147254.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@147254.4]
  input          io_DWIDTH_AXI_BID, // @[:@147254.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@147254.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@147254.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@147254.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@147254.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@147254.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@147254.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@147254.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@147254.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@147254.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@147254.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@147254.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@147254.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@147254.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@147254.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@147254.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@147254.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@147254.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@147254.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@147254.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@147254.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@147254.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@147254.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@147254.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@147254.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@147254.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@147254.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@147254.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@147254.4]
  input          io_PROTOCOL_AXI_RID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@147254.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@147254.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@147254.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@147254.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@147254.4]
  input          io_PROTOCOL_AXI_BID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@147254.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@147254.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@147254.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@147254.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@147254.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@147254.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@147254.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@147254.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@147254.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@147254.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@147254.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@147254.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@147254.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@147254.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@147254.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@147254.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@147254.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@147254.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@147254.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@147254.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@147254.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@147254.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@147254.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@147254.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@147256.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@147256.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@147256.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@147256.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@147256.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@147256.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@147256.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@147256.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@147256.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@147256.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@147398.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@147398.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@147398.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@147398.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@147398.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@147398.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@147398.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@147256.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@147398.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@147416.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@147412.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@147408.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@147407.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@147406.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@147405.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@147403.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@147402.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@147460.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@147459.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@147458.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@147457.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@147456.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@147455.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@147454.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@147453.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@147452.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@147451.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@147450.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@147448.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@147447.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@147446.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@147445.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@147444.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@147443.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@147442.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@147441.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@147440.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@147439.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@147438.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@147436.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@147435.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@147434.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@147433.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@147425.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@147420.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@147501.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@147500.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@147499.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@147498.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@147497.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@147496.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@147495.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@147494.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@147493.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@147492.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@147491.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@147489.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@147488.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@147487.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@147486.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@147485.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@147484.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@147483.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@147482.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@147481.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@147480.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@147479.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@147477.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@147476.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@147475.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@147474.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@147466.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@147461.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@147542.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@147541.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@147540.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@147539.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@147538.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@147537.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@147536.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@147535.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@147534.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@147533.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@147532.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@147530.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@147529.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@147528.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@147527.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@147526.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@147525.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@147524.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@147523.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@147522.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@147521.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@147520.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@147518.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@147517.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@147516.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@147515.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@147507.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@147502.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@147583.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@147582.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@147581.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@147580.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@147579.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@147578.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@147577.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@147576.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@147575.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@147574.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@147573.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@147571.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@147570.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@147569.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@147568.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@147567.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@147566.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@147565.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@147564.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@147563.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@147562.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@147561.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@147559.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@147558.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@147557.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@147556.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@147548.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@147543.4]
  assign accel_clock = clock; // @[:@147257.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@147258.4 Zynq.scala 54:17:@147872.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@147867.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@147860.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@147855.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@147839.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@147840.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@147841.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@147842.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@147843.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@147844.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@147845.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@147846.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@147847.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@147848.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@147849.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@147850.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@147851.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@147852.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@147853.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@147854.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@147838.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@147834.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@147829.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@147828.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@147827.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@147808.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@147792.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@147793.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@147794.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@147795.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@147796.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@147797.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@147798.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@147799.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@147800.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@147801.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@147802.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@147803.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@147804.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@147805.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@147806.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@147807.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@147791.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@147756.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@147755.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@147863.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@147862.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@147861.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@147749.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@147750.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@147753.4]
  assign FringeZynq_clock = clock; // @[:@147399.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@147400.4 Zynq.scala 53:18:@147871.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@147419.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@147418.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@147417.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@147415.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@147414.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@147413.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@147411.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@147410.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@147409.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@147404.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@147401.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@147449.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@147437.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@147432.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@147424.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@147421.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@147490.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@147478.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@147473.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@147465.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@147462.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@147531.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@147519.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@147514.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@147506.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@147503.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@147572.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@147560.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@147555.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@147547.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@147544.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@147868.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@147752.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@147751.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@147837.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@147836.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@147835.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@147833.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@147832.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@147831.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@147830.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@147866.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@147865.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@147864.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




