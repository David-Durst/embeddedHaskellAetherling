module FIFO(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  input  [7:0] I_16,
  input  [7:0] I_17,
  input  [7:0] I_18,
  input  [7:0] I_19,
  input  [7:0] I_20,
  input  [7:0] I_21,
  input  [7:0] I_22,
  input  [7:0] I_23,
  input  [7:0] I_24,
  input  [7:0] I_25,
  input  [7:0] I_26,
  input  [7:0] I_27,
  input  [7:0] I_28,
  input  [7:0] I_29,
  input  [7:0] I_30,
  input  [7:0] I_31,
  input  [7:0] I_32,
  input  [7:0] I_33,
  input  [7:0] I_34,
  input  [7:0] I_35,
  input  [7:0] I_36,
  input  [7:0] I_37,
  input  [7:0] I_38,
  input  [7:0] I_39,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15,
  output [7:0] O_16,
  output [7:0] O_17,
  output [7:0] O_18,
  output [7:0] O_19,
  output [7:0] O_20,
  output [7:0] O_21,
  output [7:0] O_22,
  output [7:0] O_23,
  output [7:0] O_24,
  output [7:0] O_25,
  output [7:0] O_26,
  output [7:0] O_27,
  output [7:0] O_28,
  output [7:0] O_29,
  output [7:0] O_30,
  output [7:0] O_31,
  output [7:0] O_32,
  output [7:0] O_33,
  output [7:0] O_34,
  output [7:0] O_35,
  output [7:0] O_36,
  output [7:0] O_37,
  output [7:0] O_38,
  output [7:0] O_39
);
  reg [7:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [7:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [7:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [7:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [7:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [7:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [7:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [7:0] _T__8; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [7:0] _T__9; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [7:0] _T__10; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [7:0] _T__11; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [7:0] _T__12; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [7:0] _T__13; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [7:0] _T__14; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [7:0] _T__15; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg [7:0] _T__16; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_16;
  reg [7:0] _T__17; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_17;
  reg [7:0] _T__18; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_18;
  reg [7:0] _T__19; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_19;
  reg [7:0] _T__20; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_20;
  reg [7:0] _T__21; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_21;
  reg [7:0] _T__22; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_22;
  reg [7:0] _T__23; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_23;
  reg [7:0] _T__24; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_24;
  reg [7:0] _T__25; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_25;
  reg [7:0] _T__26; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_26;
  reg [7:0] _T__27; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_27;
  reg [7:0] _T__28; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_28;
  reg [7:0] _T__29; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_29;
  reg [7:0] _T__30; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_30;
  reg [7:0] _T__31; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_31;
  reg [7:0] _T__32; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_32;
  reg [7:0] _T__33; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_33;
  reg [7:0] _T__34; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_34;
  reg [7:0] _T__35; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_35;
  reg [7:0] _T__36; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_36;
  reg [7:0] _T__37; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_37;
  reg [7:0] _T__38; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_38;
  reg [7:0] _T__39; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_39;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_40;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
  assign O_8 = _T__8; // @[FIFO.scala 14:7]
  assign O_9 = _T__9; // @[FIFO.scala 14:7]
  assign O_10 = _T__10; // @[FIFO.scala 14:7]
  assign O_11 = _T__11; // @[FIFO.scala 14:7]
  assign O_12 = _T__12; // @[FIFO.scala 14:7]
  assign O_13 = _T__13; // @[FIFO.scala 14:7]
  assign O_14 = _T__14; // @[FIFO.scala 14:7]
  assign O_15 = _T__15; // @[FIFO.scala 14:7]
  assign O_16 = _T__16; // @[FIFO.scala 14:7]
  assign O_17 = _T__17; // @[FIFO.scala 14:7]
  assign O_18 = _T__18; // @[FIFO.scala 14:7]
  assign O_19 = _T__19; // @[FIFO.scala 14:7]
  assign O_20 = _T__20; // @[FIFO.scala 14:7]
  assign O_21 = _T__21; // @[FIFO.scala 14:7]
  assign O_22 = _T__22; // @[FIFO.scala 14:7]
  assign O_23 = _T__23; // @[FIFO.scala 14:7]
  assign O_24 = _T__24; // @[FIFO.scala 14:7]
  assign O_25 = _T__25; // @[FIFO.scala 14:7]
  assign O_26 = _T__26; // @[FIFO.scala 14:7]
  assign O_27 = _T__27; // @[FIFO.scala 14:7]
  assign O_28 = _T__28; // @[FIFO.scala 14:7]
  assign O_29 = _T__29; // @[FIFO.scala 14:7]
  assign O_30 = _T__30; // @[FIFO.scala 14:7]
  assign O_31 = _T__31; // @[FIFO.scala 14:7]
  assign O_32 = _T__32; // @[FIFO.scala 14:7]
  assign O_33 = _T__33; // @[FIFO.scala 14:7]
  assign O_34 = _T__34; // @[FIFO.scala 14:7]
  assign O_35 = _T__35; // @[FIFO.scala 14:7]
  assign O_36 = _T__36; // @[FIFO.scala 14:7]
  assign O_37 = _T__37; // @[FIFO.scala 14:7]
  assign O_38 = _T__38; // @[FIFO.scala 14:7]
  assign O_39 = _T__39; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T__16 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T__17 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__18 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__19 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T__20 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T__21 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__22 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__23 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T__24 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T__25 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__26 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__27 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T__28 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T__29 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__30 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__31 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T__32 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T__33 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__34 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__35 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T__36 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T__37 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__38 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__39 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    _T__8 <= I_8;
    _T__9 <= I_9;
    _T__10 <= I_10;
    _T__11 <= I_11;
    _T__12 <= I_12;
    _T__13 <= I_13;
    _T__14 <= I_14;
    _T__15 <= I_15;
    _T__16 <= I_16;
    _T__17 <= I_17;
    _T__18 <= I_18;
    _T__19 <= I_19;
    _T__20 <= I_20;
    _T__21 <= I_21;
    _T__22 <= I_22;
    _T__23 <= I_23;
    _T__24 <= I_24;
    _T__25 <= I_25;
    _T__26 <= I_26;
    _T__27 <= I_27;
    _T__28 <= I_28;
    _T__29 <= I_29;
    _T__30 <= I_30;
    _T__31 <= I_31;
    _T__32 <= I_32;
    _T__33 <= I_33;
    _T__34 <= I_34;
    _T__35 <= I_35;
    _T__36 <= I_36;
    _T__37 <= I_37;
    _T__38 <= I_38;
    _T__39 <= I_39;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  output [7:0] O_t0b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
endmodule
module Add(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 108:14]
  assign O = I_t0b + 8'h5; // @[Arithmetic.scala 106:7]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n6_valid_up; // @[Top.scala 18:20]
  wire  n6_valid_down; // @[Top.scala 18:20]
  wire [7:0] n6_I0; // @[Top.scala 18:20]
  wire [7:0] n6_O_t0b; // @[Top.scala 18:20]
  wire  n7_valid_up; // @[Top.scala 22:20]
  wire  n7_valid_down; // @[Top.scala 22:20]
  wire [7:0] n7_I_t0b; // @[Top.scala 22:20]
  wire [7:0] n7_O; // @[Top.scala 22:20]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple n6 ( // @[Top.scala 18:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0(n6_I0),
    .O_t0b(n6_O_t0b)
  );
  Add n7 ( // @[Top.scala 22:20]
    .valid_up(n7_valid_up),
    .valid_down(n7_valid_down),
    .I_t0b(n7_I_t0b),
    .O(n7_O)
  );
  assign valid_down = n7_valid_down; // @[Top.scala 26:16]
  assign O = n7_O; // @[Top.scala 25:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n6_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 21:17]
  assign n6_I0 = I; // @[Top.scala 19:11]
  assign n7_valid_up = n6_valid_down; // @[Top.scala 24:17]
  assign n7_I_t0b = n6_O_t0b; // @[Top.scala 23:10]
endmodule
module MapS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  input  [7:0] I_16,
  input  [7:0] I_17,
  input  [7:0] I_18,
  input  [7:0] I_19,
  input  [7:0] I_20,
  input  [7:0] I_21,
  input  [7:0] I_22,
  input  [7:0] I_23,
  input  [7:0] I_24,
  input  [7:0] I_25,
  input  [7:0] I_26,
  input  [7:0] I_27,
  input  [7:0] I_28,
  input  [7:0] I_29,
  input  [7:0] I_30,
  input  [7:0] I_31,
  input  [7:0] I_32,
  input  [7:0] I_33,
  input  [7:0] I_34,
  input  [7:0] I_35,
  input  [7:0] I_36,
  input  [7:0] I_37,
  input  [7:0] I_38,
  input  [7:0] I_39,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15,
  output [7:0] O_16,
  output [7:0] O_17,
  output [7:0] O_18,
  output [7:0] O_19,
  output [7:0] O_20,
  output [7:0] O_21,
  output [7:0] O_22,
  output [7:0] O_23,
  output [7:0] O_24,
  output [7:0] O_25,
  output [7:0] O_26,
  output [7:0] O_27,
  output [7:0] O_28,
  output [7:0] O_29,
  output [7:0] O_30,
  output [7:0] O_31,
  output [7:0] O_32,
  output [7:0] O_33,
  output [7:0] O_34,
  output [7:0] O_35,
  output [7:0] O_36,
  output [7:0] O_37,
  output [7:0] O_38,
  output [7:0] O_39
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O; // @[MapS.scala 10:86]
  wire  other_ops_7_clock; // @[MapS.scala 10:86]
  wire  other_ops_7_reset; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O; // @[MapS.scala 10:86]
  wire  other_ops_8_clock; // @[MapS.scala 10:86]
  wire  other_ops_8_reset; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O; // @[MapS.scala 10:86]
  wire  other_ops_9_clock; // @[MapS.scala 10:86]
  wire  other_ops_9_reset; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O; // @[MapS.scala 10:86]
  wire  other_ops_10_clock; // @[MapS.scala 10:86]
  wire  other_ops_10_reset; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O; // @[MapS.scala 10:86]
  wire  other_ops_11_clock; // @[MapS.scala 10:86]
  wire  other_ops_11_reset; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O; // @[MapS.scala 10:86]
  wire  other_ops_12_clock; // @[MapS.scala 10:86]
  wire  other_ops_12_reset; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O; // @[MapS.scala 10:86]
  wire  other_ops_13_clock; // @[MapS.scala 10:86]
  wire  other_ops_13_reset; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O; // @[MapS.scala 10:86]
  wire  other_ops_14_clock; // @[MapS.scala 10:86]
  wire  other_ops_14_reset; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O; // @[MapS.scala 10:86]
  wire  other_ops_15_clock; // @[MapS.scala 10:86]
  wire  other_ops_15_reset; // @[MapS.scala 10:86]
  wire  other_ops_15_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_15_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_15_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_15_O; // @[MapS.scala 10:86]
  wire  other_ops_16_clock; // @[MapS.scala 10:86]
  wire  other_ops_16_reset; // @[MapS.scala 10:86]
  wire  other_ops_16_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_16_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_16_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_16_O; // @[MapS.scala 10:86]
  wire  other_ops_17_clock; // @[MapS.scala 10:86]
  wire  other_ops_17_reset; // @[MapS.scala 10:86]
  wire  other_ops_17_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_17_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_17_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_17_O; // @[MapS.scala 10:86]
  wire  other_ops_18_clock; // @[MapS.scala 10:86]
  wire  other_ops_18_reset; // @[MapS.scala 10:86]
  wire  other_ops_18_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_18_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_18_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_18_O; // @[MapS.scala 10:86]
  wire  other_ops_19_clock; // @[MapS.scala 10:86]
  wire  other_ops_19_reset; // @[MapS.scala 10:86]
  wire  other_ops_19_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_19_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_19_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_19_O; // @[MapS.scala 10:86]
  wire  other_ops_20_clock; // @[MapS.scala 10:86]
  wire  other_ops_20_reset; // @[MapS.scala 10:86]
  wire  other_ops_20_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_20_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_20_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_20_O; // @[MapS.scala 10:86]
  wire  other_ops_21_clock; // @[MapS.scala 10:86]
  wire  other_ops_21_reset; // @[MapS.scala 10:86]
  wire  other_ops_21_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_21_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_21_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_21_O; // @[MapS.scala 10:86]
  wire  other_ops_22_clock; // @[MapS.scala 10:86]
  wire  other_ops_22_reset; // @[MapS.scala 10:86]
  wire  other_ops_22_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_22_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_22_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_22_O; // @[MapS.scala 10:86]
  wire  other_ops_23_clock; // @[MapS.scala 10:86]
  wire  other_ops_23_reset; // @[MapS.scala 10:86]
  wire  other_ops_23_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_23_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_23_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_23_O; // @[MapS.scala 10:86]
  wire  other_ops_24_clock; // @[MapS.scala 10:86]
  wire  other_ops_24_reset; // @[MapS.scala 10:86]
  wire  other_ops_24_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_24_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_24_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_24_O; // @[MapS.scala 10:86]
  wire  other_ops_25_clock; // @[MapS.scala 10:86]
  wire  other_ops_25_reset; // @[MapS.scala 10:86]
  wire  other_ops_25_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_25_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_25_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_25_O; // @[MapS.scala 10:86]
  wire  other_ops_26_clock; // @[MapS.scala 10:86]
  wire  other_ops_26_reset; // @[MapS.scala 10:86]
  wire  other_ops_26_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_26_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_26_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_26_O; // @[MapS.scala 10:86]
  wire  other_ops_27_clock; // @[MapS.scala 10:86]
  wire  other_ops_27_reset; // @[MapS.scala 10:86]
  wire  other_ops_27_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_27_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_27_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_27_O; // @[MapS.scala 10:86]
  wire  other_ops_28_clock; // @[MapS.scala 10:86]
  wire  other_ops_28_reset; // @[MapS.scala 10:86]
  wire  other_ops_28_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_28_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_28_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_28_O; // @[MapS.scala 10:86]
  wire  other_ops_29_clock; // @[MapS.scala 10:86]
  wire  other_ops_29_reset; // @[MapS.scala 10:86]
  wire  other_ops_29_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_29_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_29_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_29_O; // @[MapS.scala 10:86]
  wire  other_ops_30_clock; // @[MapS.scala 10:86]
  wire  other_ops_30_reset; // @[MapS.scala 10:86]
  wire  other_ops_30_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_30_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_30_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_30_O; // @[MapS.scala 10:86]
  wire  other_ops_31_clock; // @[MapS.scala 10:86]
  wire  other_ops_31_reset; // @[MapS.scala 10:86]
  wire  other_ops_31_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_31_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_31_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_31_O; // @[MapS.scala 10:86]
  wire  other_ops_32_clock; // @[MapS.scala 10:86]
  wire  other_ops_32_reset; // @[MapS.scala 10:86]
  wire  other_ops_32_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_32_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_32_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_32_O; // @[MapS.scala 10:86]
  wire  other_ops_33_clock; // @[MapS.scala 10:86]
  wire  other_ops_33_reset; // @[MapS.scala 10:86]
  wire  other_ops_33_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_33_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_33_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_33_O; // @[MapS.scala 10:86]
  wire  other_ops_34_clock; // @[MapS.scala 10:86]
  wire  other_ops_34_reset; // @[MapS.scala 10:86]
  wire  other_ops_34_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_34_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_34_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_34_O; // @[MapS.scala 10:86]
  wire  other_ops_35_clock; // @[MapS.scala 10:86]
  wire  other_ops_35_reset; // @[MapS.scala 10:86]
  wire  other_ops_35_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_35_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_35_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_35_O; // @[MapS.scala 10:86]
  wire  other_ops_36_clock; // @[MapS.scala 10:86]
  wire  other_ops_36_reset; // @[MapS.scala 10:86]
  wire  other_ops_36_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_36_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_36_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_36_O; // @[MapS.scala 10:86]
  wire  other_ops_37_clock; // @[MapS.scala 10:86]
  wire  other_ops_37_reset; // @[MapS.scala 10:86]
  wire  other_ops_37_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_37_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_37_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_37_O; // @[MapS.scala 10:86]
  wire  other_ops_38_clock; // @[MapS.scala 10:86]
  wire  other_ops_38_reset; // @[MapS.scala 10:86]
  wire  other_ops_38_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_38_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_38_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_38_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  wire  _T_14; // @[MapS.scala 23:83]
  wire  _T_15; // @[MapS.scala 23:83]
  wire  _T_16; // @[MapS.scala 23:83]
  wire  _T_17; // @[MapS.scala 23:83]
  wire  _T_18; // @[MapS.scala 23:83]
  wire  _T_19; // @[MapS.scala 23:83]
  wire  _T_20; // @[MapS.scala 23:83]
  wire  _T_21; // @[MapS.scala 23:83]
  wire  _T_22; // @[MapS.scala 23:83]
  wire  _T_23; // @[MapS.scala 23:83]
  wire  _T_24; // @[MapS.scala 23:83]
  wire  _T_25; // @[MapS.scala 23:83]
  wire  _T_26; // @[MapS.scala 23:83]
  wire  _T_27; // @[MapS.scala 23:83]
  wire  _T_28; // @[MapS.scala 23:83]
  wire  _T_29; // @[MapS.scala 23:83]
  wire  _T_30; // @[MapS.scala 23:83]
  wire  _T_31; // @[MapS.scala 23:83]
  wire  _T_32; // @[MapS.scala 23:83]
  wire  _T_33; // @[MapS.scala 23:83]
  wire  _T_34; // @[MapS.scala 23:83]
  wire  _T_35; // @[MapS.scala 23:83]
  wire  _T_36; // @[MapS.scala 23:83]
  wire  _T_37; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I(other_ops_1_I),
    .O(other_ops_1_O)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I(other_ops_2_I),
    .O(other_ops_2_O)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I(other_ops_3_I),
    .O(other_ops_3_O)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I(other_ops_4_I),
    .O(other_ops_4_O)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I(other_ops_5_I),
    .O(other_ops_5_O)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I(other_ops_6_I),
    .O(other_ops_6_O)
  );
  Module_0 other_ops_7 ( // @[MapS.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I(other_ops_7_I),
    .O(other_ops_7_O)
  );
  Module_0 other_ops_8 ( // @[MapS.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I(other_ops_8_I),
    .O(other_ops_8_O)
  );
  Module_0 other_ops_9 ( // @[MapS.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I(other_ops_9_I),
    .O(other_ops_9_O)
  );
  Module_0 other_ops_10 ( // @[MapS.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I(other_ops_10_I),
    .O(other_ops_10_O)
  );
  Module_0 other_ops_11 ( // @[MapS.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I(other_ops_11_I),
    .O(other_ops_11_O)
  );
  Module_0 other_ops_12 ( // @[MapS.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I(other_ops_12_I),
    .O(other_ops_12_O)
  );
  Module_0 other_ops_13 ( // @[MapS.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I(other_ops_13_I),
    .O(other_ops_13_O)
  );
  Module_0 other_ops_14 ( // @[MapS.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I(other_ops_14_I),
    .O(other_ops_14_O)
  );
  Module_0 other_ops_15 ( // @[MapS.scala 10:86]
    .clock(other_ops_15_clock),
    .reset(other_ops_15_reset),
    .valid_up(other_ops_15_valid_up),
    .valid_down(other_ops_15_valid_down),
    .I(other_ops_15_I),
    .O(other_ops_15_O)
  );
  Module_0 other_ops_16 ( // @[MapS.scala 10:86]
    .clock(other_ops_16_clock),
    .reset(other_ops_16_reset),
    .valid_up(other_ops_16_valid_up),
    .valid_down(other_ops_16_valid_down),
    .I(other_ops_16_I),
    .O(other_ops_16_O)
  );
  Module_0 other_ops_17 ( // @[MapS.scala 10:86]
    .clock(other_ops_17_clock),
    .reset(other_ops_17_reset),
    .valid_up(other_ops_17_valid_up),
    .valid_down(other_ops_17_valid_down),
    .I(other_ops_17_I),
    .O(other_ops_17_O)
  );
  Module_0 other_ops_18 ( // @[MapS.scala 10:86]
    .clock(other_ops_18_clock),
    .reset(other_ops_18_reset),
    .valid_up(other_ops_18_valid_up),
    .valid_down(other_ops_18_valid_down),
    .I(other_ops_18_I),
    .O(other_ops_18_O)
  );
  Module_0 other_ops_19 ( // @[MapS.scala 10:86]
    .clock(other_ops_19_clock),
    .reset(other_ops_19_reset),
    .valid_up(other_ops_19_valid_up),
    .valid_down(other_ops_19_valid_down),
    .I(other_ops_19_I),
    .O(other_ops_19_O)
  );
  Module_0 other_ops_20 ( // @[MapS.scala 10:86]
    .clock(other_ops_20_clock),
    .reset(other_ops_20_reset),
    .valid_up(other_ops_20_valid_up),
    .valid_down(other_ops_20_valid_down),
    .I(other_ops_20_I),
    .O(other_ops_20_O)
  );
  Module_0 other_ops_21 ( // @[MapS.scala 10:86]
    .clock(other_ops_21_clock),
    .reset(other_ops_21_reset),
    .valid_up(other_ops_21_valid_up),
    .valid_down(other_ops_21_valid_down),
    .I(other_ops_21_I),
    .O(other_ops_21_O)
  );
  Module_0 other_ops_22 ( // @[MapS.scala 10:86]
    .clock(other_ops_22_clock),
    .reset(other_ops_22_reset),
    .valid_up(other_ops_22_valid_up),
    .valid_down(other_ops_22_valid_down),
    .I(other_ops_22_I),
    .O(other_ops_22_O)
  );
  Module_0 other_ops_23 ( // @[MapS.scala 10:86]
    .clock(other_ops_23_clock),
    .reset(other_ops_23_reset),
    .valid_up(other_ops_23_valid_up),
    .valid_down(other_ops_23_valid_down),
    .I(other_ops_23_I),
    .O(other_ops_23_O)
  );
  Module_0 other_ops_24 ( // @[MapS.scala 10:86]
    .clock(other_ops_24_clock),
    .reset(other_ops_24_reset),
    .valid_up(other_ops_24_valid_up),
    .valid_down(other_ops_24_valid_down),
    .I(other_ops_24_I),
    .O(other_ops_24_O)
  );
  Module_0 other_ops_25 ( // @[MapS.scala 10:86]
    .clock(other_ops_25_clock),
    .reset(other_ops_25_reset),
    .valid_up(other_ops_25_valid_up),
    .valid_down(other_ops_25_valid_down),
    .I(other_ops_25_I),
    .O(other_ops_25_O)
  );
  Module_0 other_ops_26 ( // @[MapS.scala 10:86]
    .clock(other_ops_26_clock),
    .reset(other_ops_26_reset),
    .valid_up(other_ops_26_valid_up),
    .valid_down(other_ops_26_valid_down),
    .I(other_ops_26_I),
    .O(other_ops_26_O)
  );
  Module_0 other_ops_27 ( // @[MapS.scala 10:86]
    .clock(other_ops_27_clock),
    .reset(other_ops_27_reset),
    .valid_up(other_ops_27_valid_up),
    .valid_down(other_ops_27_valid_down),
    .I(other_ops_27_I),
    .O(other_ops_27_O)
  );
  Module_0 other_ops_28 ( // @[MapS.scala 10:86]
    .clock(other_ops_28_clock),
    .reset(other_ops_28_reset),
    .valid_up(other_ops_28_valid_up),
    .valid_down(other_ops_28_valid_down),
    .I(other_ops_28_I),
    .O(other_ops_28_O)
  );
  Module_0 other_ops_29 ( // @[MapS.scala 10:86]
    .clock(other_ops_29_clock),
    .reset(other_ops_29_reset),
    .valid_up(other_ops_29_valid_up),
    .valid_down(other_ops_29_valid_down),
    .I(other_ops_29_I),
    .O(other_ops_29_O)
  );
  Module_0 other_ops_30 ( // @[MapS.scala 10:86]
    .clock(other_ops_30_clock),
    .reset(other_ops_30_reset),
    .valid_up(other_ops_30_valid_up),
    .valid_down(other_ops_30_valid_down),
    .I(other_ops_30_I),
    .O(other_ops_30_O)
  );
  Module_0 other_ops_31 ( // @[MapS.scala 10:86]
    .clock(other_ops_31_clock),
    .reset(other_ops_31_reset),
    .valid_up(other_ops_31_valid_up),
    .valid_down(other_ops_31_valid_down),
    .I(other_ops_31_I),
    .O(other_ops_31_O)
  );
  Module_0 other_ops_32 ( // @[MapS.scala 10:86]
    .clock(other_ops_32_clock),
    .reset(other_ops_32_reset),
    .valid_up(other_ops_32_valid_up),
    .valid_down(other_ops_32_valid_down),
    .I(other_ops_32_I),
    .O(other_ops_32_O)
  );
  Module_0 other_ops_33 ( // @[MapS.scala 10:86]
    .clock(other_ops_33_clock),
    .reset(other_ops_33_reset),
    .valid_up(other_ops_33_valid_up),
    .valid_down(other_ops_33_valid_down),
    .I(other_ops_33_I),
    .O(other_ops_33_O)
  );
  Module_0 other_ops_34 ( // @[MapS.scala 10:86]
    .clock(other_ops_34_clock),
    .reset(other_ops_34_reset),
    .valid_up(other_ops_34_valid_up),
    .valid_down(other_ops_34_valid_down),
    .I(other_ops_34_I),
    .O(other_ops_34_O)
  );
  Module_0 other_ops_35 ( // @[MapS.scala 10:86]
    .clock(other_ops_35_clock),
    .reset(other_ops_35_reset),
    .valid_up(other_ops_35_valid_up),
    .valid_down(other_ops_35_valid_down),
    .I(other_ops_35_I),
    .O(other_ops_35_O)
  );
  Module_0 other_ops_36 ( // @[MapS.scala 10:86]
    .clock(other_ops_36_clock),
    .reset(other_ops_36_reset),
    .valid_up(other_ops_36_valid_up),
    .valid_down(other_ops_36_valid_down),
    .I(other_ops_36_I),
    .O(other_ops_36_O)
  );
  Module_0 other_ops_37 ( // @[MapS.scala 10:86]
    .clock(other_ops_37_clock),
    .reset(other_ops_37_reset),
    .valid_up(other_ops_37_valid_up),
    .valid_down(other_ops_37_valid_down),
    .I(other_ops_37_I),
    .O(other_ops_37_O)
  );
  Module_0 other_ops_38 ( // @[MapS.scala 10:86]
    .clock(other_ops_38_clock),
    .reset(other_ops_38_reset),
    .valid_up(other_ops_38_valid_up),
    .valid_down(other_ops_38_valid_down),
    .I(other_ops_38_I),
    .O(other_ops_38_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign _T_14 = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:83]
  assign _T_15 = _T_14 & other_ops_15_valid_down; // @[MapS.scala 23:83]
  assign _T_16 = _T_15 & other_ops_16_valid_down; // @[MapS.scala 23:83]
  assign _T_17 = _T_16 & other_ops_17_valid_down; // @[MapS.scala 23:83]
  assign _T_18 = _T_17 & other_ops_18_valid_down; // @[MapS.scala 23:83]
  assign _T_19 = _T_18 & other_ops_19_valid_down; // @[MapS.scala 23:83]
  assign _T_20 = _T_19 & other_ops_20_valid_down; // @[MapS.scala 23:83]
  assign _T_21 = _T_20 & other_ops_21_valid_down; // @[MapS.scala 23:83]
  assign _T_22 = _T_21 & other_ops_22_valid_down; // @[MapS.scala 23:83]
  assign _T_23 = _T_22 & other_ops_23_valid_down; // @[MapS.scala 23:83]
  assign _T_24 = _T_23 & other_ops_24_valid_down; // @[MapS.scala 23:83]
  assign _T_25 = _T_24 & other_ops_25_valid_down; // @[MapS.scala 23:83]
  assign _T_26 = _T_25 & other_ops_26_valid_down; // @[MapS.scala 23:83]
  assign _T_27 = _T_26 & other_ops_27_valid_down; // @[MapS.scala 23:83]
  assign _T_28 = _T_27 & other_ops_28_valid_down; // @[MapS.scala 23:83]
  assign _T_29 = _T_28 & other_ops_29_valid_down; // @[MapS.scala 23:83]
  assign _T_30 = _T_29 & other_ops_30_valid_down; // @[MapS.scala 23:83]
  assign _T_31 = _T_30 & other_ops_31_valid_down; // @[MapS.scala 23:83]
  assign _T_32 = _T_31 & other_ops_32_valid_down; // @[MapS.scala 23:83]
  assign _T_33 = _T_32 & other_ops_33_valid_down; // @[MapS.scala 23:83]
  assign _T_34 = _T_33 & other_ops_34_valid_down; // @[MapS.scala 23:83]
  assign _T_35 = _T_34 & other_ops_35_valid_down; // @[MapS.scala 23:83]
  assign _T_36 = _T_35 & other_ops_36_valid_down; // @[MapS.scala 23:83]
  assign _T_37 = _T_36 & other_ops_37_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_37 & other_ops_38_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign O_8 = other_ops_7_O; // @[MapS.scala 21:12]
  assign O_9 = other_ops_8_O; // @[MapS.scala 21:12]
  assign O_10 = other_ops_9_O; // @[MapS.scala 21:12]
  assign O_11 = other_ops_10_O; // @[MapS.scala 21:12]
  assign O_12 = other_ops_11_O; // @[MapS.scala 21:12]
  assign O_13 = other_ops_12_O; // @[MapS.scala 21:12]
  assign O_14 = other_ops_13_O; // @[MapS.scala 21:12]
  assign O_15 = other_ops_14_O; // @[MapS.scala 21:12]
  assign O_16 = other_ops_15_O; // @[MapS.scala 21:12]
  assign O_17 = other_ops_16_O; // @[MapS.scala 21:12]
  assign O_18 = other_ops_17_O; // @[MapS.scala 21:12]
  assign O_19 = other_ops_18_O; // @[MapS.scala 21:12]
  assign O_20 = other_ops_19_O; // @[MapS.scala 21:12]
  assign O_21 = other_ops_20_O; // @[MapS.scala 21:12]
  assign O_22 = other_ops_21_O; // @[MapS.scala 21:12]
  assign O_23 = other_ops_22_O; // @[MapS.scala 21:12]
  assign O_24 = other_ops_23_O; // @[MapS.scala 21:12]
  assign O_25 = other_ops_24_O; // @[MapS.scala 21:12]
  assign O_26 = other_ops_25_O; // @[MapS.scala 21:12]
  assign O_27 = other_ops_26_O; // @[MapS.scala 21:12]
  assign O_28 = other_ops_27_O; // @[MapS.scala 21:12]
  assign O_29 = other_ops_28_O; // @[MapS.scala 21:12]
  assign O_30 = other_ops_29_O; // @[MapS.scala 21:12]
  assign O_31 = other_ops_30_O; // @[MapS.scala 21:12]
  assign O_32 = other_ops_31_O; // @[MapS.scala 21:12]
  assign O_33 = other_ops_32_O; // @[MapS.scala 21:12]
  assign O_34 = other_ops_33_O; // @[MapS.scala 21:12]
  assign O_35 = other_ops_34_O; // @[MapS.scala 21:12]
  assign O_36 = other_ops_35_O; // @[MapS.scala 21:12]
  assign O_37 = other_ops_36_O; // @[MapS.scala 21:12]
  assign O_38 = other_ops_37_O; // @[MapS.scala 21:12]
  assign O_39 = other_ops_38_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I = I_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I = I_3; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I = I_4; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I = I_5; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I = I_6; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I = I_7; // @[MapS.scala 20:41]
  assign other_ops_7_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_7_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I = I_8; // @[MapS.scala 20:41]
  assign other_ops_8_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_8_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I = I_9; // @[MapS.scala 20:41]
  assign other_ops_9_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_9_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I = I_10; // @[MapS.scala 20:41]
  assign other_ops_10_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_10_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I = I_11; // @[MapS.scala 20:41]
  assign other_ops_11_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_11_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I = I_12; // @[MapS.scala 20:41]
  assign other_ops_12_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_12_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I = I_13; // @[MapS.scala 20:41]
  assign other_ops_13_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_13_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I = I_14; // @[MapS.scala 20:41]
  assign other_ops_14_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_14_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I = I_15; // @[MapS.scala 20:41]
  assign other_ops_15_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_15_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_15_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_15_I = I_16; // @[MapS.scala 20:41]
  assign other_ops_16_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_16_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_16_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_16_I = I_17; // @[MapS.scala 20:41]
  assign other_ops_17_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_17_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_17_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_17_I = I_18; // @[MapS.scala 20:41]
  assign other_ops_18_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_18_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_18_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_18_I = I_19; // @[MapS.scala 20:41]
  assign other_ops_19_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_19_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_19_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_19_I = I_20; // @[MapS.scala 20:41]
  assign other_ops_20_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_20_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_20_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_20_I = I_21; // @[MapS.scala 20:41]
  assign other_ops_21_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_21_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_21_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_21_I = I_22; // @[MapS.scala 20:41]
  assign other_ops_22_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_22_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_22_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_22_I = I_23; // @[MapS.scala 20:41]
  assign other_ops_23_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_23_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_23_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_23_I = I_24; // @[MapS.scala 20:41]
  assign other_ops_24_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_24_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_24_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_24_I = I_25; // @[MapS.scala 20:41]
  assign other_ops_25_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_25_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_25_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_25_I = I_26; // @[MapS.scala 20:41]
  assign other_ops_26_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_26_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_26_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_26_I = I_27; // @[MapS.scala 20:41]
  assign other_ops_27_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_27_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_27_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_27_I = I_28; // @[MapS.scala 20:41]
  assign other_ops_28_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_28_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_28_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_28_I = I_29; // @[MapS.scala 20:41]
  assign other_ops_29_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_29_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_29_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_29_I = I_30; // @[MapS.scala 20:41]
  assign other_ops_30_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_30_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_30_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_30_I = I_31; // @[MapS.scala 20:41]
  assign other_ops_31_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_31_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_31_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_31_I = I_32; // @[MapS.scala 20:41]
  assign other_ops_32_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_32_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_32_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_32_I = I_33; // @[MapS.scala 20:41]
  assign other_ops_33_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_33_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_33_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_33_I = I_34; // @[MapS.scala 20:41]
  assign other_ops_34_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_34_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_34_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_34_I = I_35; // @[MapS.scala 20:41]
  assign other_ops_35_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_35_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_35_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_35_I = I_36; // @[MapS.scala 20:41]
  assign other_ops_36_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_36_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_36_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_36_I = I_37; // @[MapS.scala 20:41]
  assign other_ops_37_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_37_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_37_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_37_I = I_38; // @[MapS.scala 20:41]
  assign other_ops_38_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_38_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_38_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_38_I = I_39; // @[MapS.scala 20:41]
endmodule
module MapT(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  input  [7:0] I_16,
  input  [7:0] I_17,
  input  [7:0] I_18,
  input  [7:0] I_19,
  input  [7:0] I_20,
  input  [7:0] I_21,
  input  [7:0] I_22,
  input  [7:0] I_23,
  input  [7:0] I_24,
  input  [7:0] I_25,
  input  [7:0] I_26,
  input  [7:0] I_27,
  input  [7:0] I_28,
  input  [7:0] I_29,
  input  [7:0] I_30,
  input  [7:0] I_31,
  input  [7:0] I_32,
  input  [7:0] I_33,
  input  [7:0] I_34,
  input  [7:0] I_35,
  input  [7:0] I_36,
  input  [7:0] I_37,
  input  [7:0] I_38,
  input  [7:0] I_39,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15,
  output [7:0] O_16,
  output [7:0] O_17,
  output [7:0] O_18,
  output [7:0] O_19,
  output [7:0] O_20,
  output [7:0] O_21,
  output [7:0] O_22,
  output [7:0] O_23,
  output [7:0] O_24,
  output [7:0] O_25,
  output [7:0] O_26,
  output [7:0] O_27,
  output [7:0] O_28,
  output [7:0] O_29,
  output [7:0] O_30,
  output [7:0] O_31,
  output [7:0] O_32,
  output [7:0] O_33,
  output [7:0] O_34,
  output [7:0] O_35,
  output [7:0] O_36,
  output [7:0] O_37,
  output [7:0] O_38,
  output [7:0] O_39
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3; // @[MapT.scala 8:20]
  wire [7:0] op_I_4; // @[MapT.scala 8:20]
  wire [7:0] op_I_5; // @[MapT.scala 8:20]
  wire [7:0] op_I_6; // @[MapT.scala 8:20]
  wire [7:0] op_I_7; // @[MapT.scala 8:20]
  wire [7:0] op_I_8; // @[MapT.scala 8:20]
  wire [7:0] op_I_9; // @[MapT.scala 8:20]
  wire [7:0] op_I_10; // @[MapT.scala 8:20]
  wire [7:0] op_I_11; // @[MapT.scala 8:20]
  wire [7:0] op_I_12; // @[MapT.scala 8:20]
  wire [7:0] op_I_13; // @[MapT.scala 8:20]
  wire [7:0] op_I_14; // @[MapT.scala 8:20]
  wire [7:0] op_I_15; // @[MapT.scala 8:20]
  wire [7:0] op_I_16; // @[MapT.scala 8:20]
  wire [7:0] op_I_17; // @[MapT.scala 8:20]
  wire [7:0] op_I_18; // @[MapT.scala 8:20]
  wire [7:0] op_I_19; // @[MapT.scala 8:20]
  wire [7:0] op_I_20; // @[MapT.scala 8:20]
  wire [7:0] op_I_21; // @[MapT.scala 8:20]
  wire [7:0] op_I_22; // @[MapT.scala 8:20]
  wire [7:0] op_I_23; // @[MapT.scala 8:20]
  wire [7:0] op_I_24; // @[MapT.scala 8:20]
  wire [7:0] op_I_25; // @[MapT.scala 8:20]
  wire [7:0] op_I_26; // @[MapT.scala 8:20]
  wire [7:0] op_I_27; // @[MapT.scala 8:20]
  wire [7:0] op_I_28; // @[MapT.scala 8:20]
  wire [7:0] op_I_29; // @[MapT.scala 8:20]
  wire [7:0] op_I_30; // @[MapT.scala 8:20]
  wire [7:0] op_I_31; // @[MapT.scala 8:20]
  wire [7:0] op_I_32; // @[MapT.scala 8:20]
  wire [7:0] op_I_33; // @[MapT.scala 8:20]
  wire [7:0] op_I_34; // @[MapT.scala 8:20]
  wire [7:0] op_I_35; // @[MapT.scala 8:20]
  wire [7:0] op_I_36; // @[MapT.scala 8:20]
  wire [7:0] op_I_37; // @[MapT.scala 8:20]
  wire [7:0] op_I_38; // @[MapT.scala 8:20]
  wire [7:0] op_I_39; // @[MapT.scala 8:20]
  wire [7:0] op_O_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3; // @[MapT.scala 8:20]
  wire [7:0] op_O_4; // @[MapT.scala 8:20]
  wire [7:0] op_O_5; // @[MapT.scala 8:20]
  wire [7:0] op_O_6; // @[MapT.scala 8:20]
  wire [7:0] op_O_7; // @[MapT.scala 8:20]
  wire [7:0] op_O_8; // @[MapT.scala 8:20]
  wire [7:0] op_O_9; // @[MapT.scala 8:20]
  wire [7:0] op_O_10; // @[MapT.scala 8:20]
  wire [7:0] op_O_11; // @[MapT.scala 8:20]
  wire [7:0] op_O_12; // @[MapT.scala 8:20]
  wire [7:0] op_O_13; // @[MapT.scala 8:20]
  wire [7:0] op_O_14; // @[MapT.scala 8:20]
  wire [7:0] op_O_15; // @[MapT.scala 8:20]
  wire [7:0] op_O_16; // @[MapT.scala 8:20]
  wire [7:0] op_O_17; // @[MapT.scala 8:20]
  wire [7:0] op_O_18; // @[MapT.scala 8:20]
  wire [7:0] op_O_19; // @[MapT.scala 8:20]
  wire [7:0] op_O_20; // @[MapT.scala 8:20]
  wire [7:0] op_O_21; // @[MapT.scala 8:20]
  wire [7:0] op_O_22; // @[MapT.scala 8:20]
  wire [7:0] op_O_23; // @[MapT.scala 8:20]
  wire [7:0] op_O_24; // @[MapT.scala 8:20]
  wire [7:0] op_O_25; // @[MapT.scala 8:20]
  wire [7:0] op_O_26; // @[MapT.scala 8:20]
  wire [7:0] op_O_27; // @[MapT.scala 8:20]
  wire [7:0] op_O_28; // @[MapT.scala 8:20]
  wire [7:0] op_O_29; // @[MapT.scala 8:20]
  wire [7:0] op_O_30; // @[MapT.scala 8:20]
  wire [7:0] op_O_31; // @[MapT.scala 8:20]
  wire [7:0] op_O_32; // @[MapT.scala 8:20]
  wire [7:0] op_O_33; // @[MapT.scala 8:20]
  wire [7:0] op_O_34; // @[MapT.scala 8:20]
  wire [7:0] op_O_35; // @[MapT.scala 8:20]
  wire [7:0] op_O_36; // @[MapT.scala 8:20]
  wire [7:0] op_O_37; // @[MapT.scala 8:20]
  wire [7:0] op_O_38; // @[MapT.scala 8:20]
  wire [7:0] op_O_39; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .I_3(op_I_3),
    .I_4(op_I_4),
    .I_5(op_I_5),
    .I_6(op_I_6),
    .I_7(op_I_7),
    .I_8(op_I_8),
    .I_9(op_I_9),
    .I_10(op_I_10),
    .I_11(op_I_11),
    .I_12(op_I_12),
    .I_13(op_I_13),
    .I_14(op_I_14),
    .I_15(op_I_15),
    .I_16(op_I_16),
    .I_17(op_I_17),
    .I_18(op_I_18),
    .I_19(op_I_19),
    .I_20(op_I_20),
    .I_21(op_I_21),
    .I_22(op_I_22),
    .I_23(op_I_23),
    .I_24(op_I_24),
    .I_25(op_I_25),
    .I_26(op_I_26),
    .I_27(op_I_27),
    .I_28(op_I_28),
    .I_29(op_I_29),
    .I_30(op_I_30),
    .I_31(op_I_31),
    .I_32(op_I_32),
    .I_33(op_I_33),
    .I_34(op_I_34),
    .I_35(op_I_35),
    .I_36(op_I_36),
    .I_37(op_I_37),
    .I_38(op_I_38),
    .I_39(op_I_39),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7),
    .O_8(op_O_8),
    .O_9(op_O_9),
    .O_10(op_O_10),
    .O_11(op_O_11),
    .O_12(op_O_12),
    .O_13(op_O_13),
    .O_14(op_O_14),
    .O_15(op_O_15),
    .O_16(op_O_16),
    .O_17(op_O_17),
    .O_18(op_O_18),
    .O_19(op_O_19),
    .O_20(op_O_20),
    .O_21(op_O_21),
    .O_22(op_O_22),
    .O_23(op_O_23),
    .O_24(op_O_24),
    .O_25(op_O_25),
    .O_26(op_O_26),
    .O_27(op_O_27),
    .O_28(op_O_28),
    .O_29(op_O_29),
    .O_30(op_O_30),
    .O_31(op_O_31),
    .O_32(op_O_32),
    .O_33(op_O_33),
    .O_34(op_O_34),
    .O_35(op_O_35),
    .O_36(op_O_36),
    .O_37(op_O_37),
    .O_38(op_O_38),
    .O_39(op_O_39)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign O_8 = op_O_8; // @[MapT.scala 15:7]
  assign O_9 = op_O_9; // @[MapT.scala 15:7]
  assign O_10 = op_O_10; // @[MapT.scala 15:7]
  assign O_11 = op_O_11; // @[MapT.scala 15:7]
  assign O_12 = op_O_12; // @[MapT.scala 15:7]
  assign O_13 = op_O_13; // @[MapT.scala 15:7]
  assign O_14 = op_O_14; // @[MapT.scala 15:7]
  assign O_15 = op_O_15; // @[MapT.scala 15:7]
  assign O_16 = op_O_16; // @[MapT.scala 15:7]
  assign O_17 = op_O_17; // @[MapT.scala 15:7]
  assign O_18 = op_O_18; // @[MapT.scala 15:7]
  assign O_19 = op_O_19; // @[MapT.scala 15:7]
  assign O_20 = op_O_20; // @[MapT.scala 15:7]
  assign O_21 = op_O_21; // @[MapT.scala 15:7]
  assign O_22 = op_O_22; // @[MapT.scala 15:7]
  assign O_23 = op_O_23; // @[MapT.scala 15:7]
  assign O_24 = op_O_24; // @[MapT.scala 15:7]
  assign O_25 = op_O_25; // @[MapT.scala 15:7]
  assign O_26 = op_O_26; // @[MapT.scala 15:7]
  assign O_27 = op_O_27; // @[MapT.scala 15:7]
  assign O_28 = op_O_28; // @[MapT.scala 15:7]
  assign O_29 = op_O_29; // @[MapT.scala 15:7]
  assign O_30 = op_O_30; // @[MapT.scala 15:7]
  assign O_31 = op_O_31; // @[MapT.scala 15:7]
  assign O_32 = op_O_32; // @[MapT.scala 15:7]
  assign O_33 = op_O_33; // @[MapT.scala 15:7]
  assign O_34 = op_O_34; // @[MapT.scala 15:7]
  assign O_35 = op_O_35; // @[MapT.scala 15:7]
  assign O_36 = op_O_36; // @[MapT.scala 15:7]
  assign O_37 = op_O_37; // @[MapT.scala 15:7]
  assign O_38 = op_O_38; // @[MapT.scala 15:7]
  assign O_39 = op_O_39; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
  assign op_I_3 = I_3; // @[MapT.scala 14:10]
  assign op_I_4 = I_4; // @[MapT.scala 14:10]
  assign op_I_5 = I_5; // @[MapT.scala 14:10]
  assign op_I_6 = I_6; // @[MapT.scala 14:10]
  assign op_I_7 = I_7; // @[MapT.scala 14:10]
  assign op_I_8 = I_8; // @[MapT.scala 14:10]
  assign op_I_9 = I_9; // @[MapT.scala 14:10]
  assign op_I_10 = I_10; // @[MapT.scala 14:10]
  assign op_I_11 = I_11; // @[MapT.scala 14:10]
  assign op_I_12 = I_12; // @[MapT.scala 14:10]
  assign op_I_13 = I_13; // @[MapT.scala 14:10]
  assign op_I_14 = I_14; // @[MapT.scala 14:10]
  assign op_I_15 = I_15; // @[MapT.scala 14:10]
  assign op_I_16 = I_16; // @[MapT.scala 14:10]
  assign op_I_17 = I_17; // @[MapT.scala 14:10]
  assign op_I_18 = I_18; // @[MapT.scala 14:10]
  assign op_I_19 = I_19; // @[MapT.scala 14:10]
  assign op_I_20 = I_20; // @[MapT.scala 14:10]
  assign op_I_21 = I_21; // @[MapT.scala 14:10]
  assign op_I_22 = I_22; // @[MapT.scala 14:10]
  assign op_I_23 = I_23; // @[MapT.scala 14:10]
  assign op_I_24 = I_24; // @[MapT.scala 14:10]
  assign op_I_25 = I_25; // @[MapT.scala 14:10]
  assign op_I_26 = I_26; // @[MapT.scala 14:10]
  assign op_I_27 = I_27; // @[MapT.scala 14:10]
  assign op_I_28 = I_28; // @[MapT.scala 14:10]
  assign op_I_29 = I_29; // @[MapT.scala 14:10]
  assign op_I_30 = I_30; // @[MapT.scala 14:10]
  assign op_I_31 = I_31; // @[MapT.scala 14:10]
  assign op_I_32 = I_32; // @[MapT.scala 14:10]
  assign op_I_33 = I_33; // @[MapT.scala 14:10]
  assign op_I_34 = I_34; // @[MapT.scala 14:10]
  assign op_I_35 = I_35; // @[MapT.scala 14:10]
  assign op_I_36 = I_36; // @[MapT.scala 14:10]
  assign op_I_37 = I_37; // @[MapT.scala 14:10]
  assign op_I_38 = I_38; // @[MapT.scala 14:10]
  assign op_I_39 = I_39; // @[MapT.scala 14:10]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  input  [7:0] I_16,
  input  [7:0] I_17,
  input  [7:0] I_18,
  input  [7:0] I_19,
  input  [7:0] I_20,
  input  [7:0] I_21,
  input  [7:0] I_22,
  input  [7:0] I_23,
  input  [7:0] I_24,
  input  [7:0] I_25,
  input  [7:0] I_26,
  input  [7:0] I_27,
  input  [7:0] I_28,
  input  [7:0] I_29,
  input  [7:0] I_30,
  input  [7:0] I_31,
  input  [7:0] I_32,
  input  [7:0] I_33,
  input  [7:0] I_34,
  input  [7:0] I_35,
  input  [7:0] I_36,
  input  [7:0] I_37,
  input  [7:0] I_38,
  input  [7:0] I_39,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15,
  output [7:0] O_16,
  output [7:0] O_17,
  output [7:0] O_18,
  output [7:0] O_19,
  output [7:0] O_20,
  output [7:0] O_21,
  output [7:0] O_22,
  output [7:0] O_23,
  output [7:0] O_24,
  output [7:0] O_25,
  output [7:0] O_26,
  output [7:0] O_27,
  output [7:0] O_28,
  output [7:0] O_29,
  output [7:0] O_30,
  output [7:0] O_31,
  output [7:0] O_32,
  output [7:0] O_33,
  output [7:0] O_34,
  output [7:0] O_35,
  output [7:0] O_36,
  output [7:0] O_37,
  output [7:0] O_38,
  output [7:0] O_39
);
  wire  n1_clock; // @[Top.scala 32:20]
  wire  n1_reset; // @[Top.scala 32:20]
  wire  n1_valid_up; // @[Top.scala 32:20]
  wire  n1_valid_down; // @[Top.scala 32:20]
  wire [7:0] n1_I_0; // @[Top.scala 32:20]
  wire [7:0] n1_I_1; // @[Top.scala 32:20]
  wire [7:0] n1_I_2; // @[Top.scala 32:20]
  wire [7:0] n1_I_3; // @[Top.scala 32:20]
  wire [7:0] n1_I_4; // @[Top.scala 32:20]
  wire [7:0] n1_I_5; // @[Top.scala 32:20]
  wire [7:0] n1_I_6; // @[Top.scala 32:20]
  wire [7:0] n1_I_7; // @[Top.scala 32:20]
  wire [7:0] n1_I_8; // @[Top.scala 32:20]
  wire [7:0] n1_I_9; // @[Top.scala 32:20]
  wire [7:0] n1_I_10; // @[Top.scala 32:20]
  wire [7:0] n1_I_11; // @[Top.scala 32:20]
  wire [7:0] n1_I_12; // @[Top.scala 32:20]
  wire [7:0] n1_I_13; // @[Top.scala 32:20]
  wire [7:0] n1_I_14; // @[Top.scala 32:20]
  wire [7:0] n1_I_15; // @[Top.scala 32:20]
  wire [7:0] n1_I_16; // @[Top.scala 32:20]
  wire [7:0] n1_I_17; // @[Top.scala 32:20]
  wire [7:0] n1_I_18; // @[Top.scala 32:20]
  wire [7:0] n1_I_19; // @[Top.scala 32:20]
  wire [7:0] n1_I_20; // @[Top.scala 32:20]
  wire [7:0] n1_I_21; // @[Top.scala 32:20]
  wire [7:0] n1_I_22; // @[Top.scala 32:20]
  wire [7:0] n1_I_23; // @[Top.scala 32:20]
  wire [7:0] n1_I_24; // @[Top.scala 32:20]
  wire [7:0] n1_I_25; // @[Top.scala 32:20]
  wire [7:0] n1_I_26; // @[Top.scala 32:20]
  wire [7:0] n1_I_27; // @[Top.scala 32:20]
  wire [7:0] n1_I_28; // @[Top.scala 32:20]
  wire [7:0] n1_I_29; // @[Top.scala 32:20]
  wire [7:0] n1_I_30; // @[Top.scala 32:20]
  wire [7:0] n1_I_31; // @[Top.scala 32:20]
  wire [7:0] n1_I_32; // @[Top.scala 32:20]
  wire [7:0] n1_I_33; // @[Top.scala 32:20]
  wire [7:0] n1_I_34; // @[Top.scala 32:20]
  wire [7:0] n1_I_35; // @[Top.scala 32:20]
  wire [7:0] n1_I_36; // @[Top.scala 32:20]
  wire [7:0] n1_I_37; // @[Top.scala 32:20]
  wire [7:0] n1_I_38; // @[Top.scala 32:20]
  wire [7:0] n1_I_39; // @[Top.scala 32:20]
  wire [7:0] n1_O_0; // @[Top.scala 32:20]
  wire [7:0] n1_O_1; // @[Top.scala 32:20]
  wire [7:0] n1_O_2; // @[Top.scala 32:20]
  wire [7:0] n1_O_3; // @[Top.scala 32:20]
  wire [7:0] n1_O_4; // @[Top.scala 32:20]
  wire [7:0] n1_O_5; // @[Top.scala 32:20]
  wire [7:0] n1_O_6; // @[Top.scala 32:20]
  wire [7:0] n1_O_7; // @[Top.scala 32:20]
  wire [7:0] n1_O_8; // @[Top.scala 32:20]
  wire [7:0] n1_O_9; // @[Top.scala 32:20]
  wire [7:0] n1_O_10; // @[Top.scala 32:20]
  wire [7:0] n1_O_11; // @[Top.scala 32:20]
  wire [7:0] n1_O_12; // @[Top.scala 32:20]
  wire [7:0] n1_O_13; // @[Top.scala 32:20]
  wire [7:0] n1_O_14; // @[Top.scala 32:20]
  wire [7:0] n1_O_15; // @[Top.scala 32:20]
  wire [7:0] n1_O_16; // @[Top.scala 32:20]
  wire [7:0] n1_O_17; // @[Top.scala 32:20]
  wire [7:0] n1_O_18; // @[Top.scala 32:20]
  wire [7:0] n1_O_19; // @[Top.scala 32:20]
  wire [7:0] n1_O_20; // @[Top.scala 32:20]
  wire [7:0] n1_O_21; // @[Top.scala 32:20]
  wire [7:0] n1_O_22; // @[Top.scala 32:20]
  wire [7:0] n1_O_23; // @[Top.scala 32:20]
  wire [7:0] n1_O_24; // @[Top.scala 32:20]
  wire [7:0] n1_O_25; // @[Top.scala 32:20]
  wire [7:0] n1_O_26; // @[Top.scala 32:20]
  wire [7:0] n1_O_27; // @[Top.scala 32:20]
  wire [7:0] n1_O_28; // @[Top.scala 32:20]
  wire [7:0] n1_O_29; // @[Top.scala 32:20]
  wire [7:0] n1_O_30; // @[Top.scala 32:20]
  wire [7:0] n1_O_31; // @[Top.scala 32:20]
  wire [7:0] n1_O_32; // @[Top.scala 32:20]
  wire [7:0] n1_O_33; // @[Top.scala 32:20]
  wire [7:0] n1_O_34; // @[Top.scala 32:20]
  wire [7:0] n1_O_35; // @[Top.scala 32:20]
  wire [7:0] n1_O_36; // @[Top.scala 32:20]
  wire [7:0] n1_O_37; // @[Top.scala 32:20]
  wire [7:0] n1_O_38; // @[Top.scala 32:20]
  wire [7:0] n1_O_39; // @[Top.scala 32:20]
  wire  n9_clock; // @[Top.scala 35:20]
  wire  n9_reset; // @[Top.scala 35:20]
  wire  n9_valid_up; // @[Top.scala 35:20]
  wire  n9_valid_down; // @[Top.scala 35:20]
  wire [7:0] n9_I_0; // @[Top.scala 35:20]
  wire [7:0] n9_I_1; // @[Top.scala 35:20]
  wire [7:0] n9_I_2; // @[Top.scala 35:20]
  wire [7:0] n9_I_3; // @[Top.scala 35:20]
  wire [7:0] n9_I_4; // @[Top.scala 35:20]
  wire [7:0] n9_I_5; // @[Top.scala 35:20]
  wire [7:0] n9_I_6; // @[Top.scala 35:20]
  wire [7:0] n9_I_7; // @[Top.scala 35:20]
  wire [7:0] n9_I_8; // @[Top.scala 35:20]
  wire [7:0] n9_I_9; // @[Top.scala 35:20]
  wire [7:0] n9_I_10; // @[Top.scala 35:20]
  wire [7:0] n9_I_11; // @[Top.scala 35:20]
  wire [7:0] n9_I_12; // @[Top.scala 35:20]
  wire [7:0] n9_I_13; // @[Top.scala 35:20]
  wire [7:0] n9_I_14; // @[Top.scala 35:20]
  wire [7:0] n9_I_15; // @[Top.scala 35:20]
  wire [7:0] n9_I_16; // @[Top.scala 35:20]
  wire [7:0] n9_I_17; // @[Top.scala 35:20]
  wire [7:0] n9_I_18; // @[Top.scala 35:20]
  wire [7:0] n9_I_19; // @[Top.scala 35:20]
  wire [7:0] n9_I_20; // @[Top.scala 35:20]
  wire [7:0] n9_I_21; // @[Top.scala 35:20]
  wire [7:0] n9_I_22; // @[Top.scala 35:20]
  wire [7:0] n9_I_23; // @[Top.scala 35:20]
  wire [7:0] n9_I_24; // @[Top.scala 35:20]
  wire [7:0] n9_I_25; // @[Top.scala 35:20]
  wire [7:0] n9_I_26; // @[Top.scala 35:20]
  wire [7:0] n9_I_27; // @[Top.scala 35:20]
  wire [7:0] n9_I_28; // @[Top.scala 35:20]
  wire [7:0] n9_I_29; // @[Top.scala 35:20]
  wire [7:0] n9_I_30; // @[Top.scala 35:20]
  wire [7:0] n9_I_31; // @[Top.scala 35:20]
  wire [7:0] n9_I_32; // @[Top.scala 35:20]
  wire [7:0] n9_I_33; // @[Top.scala 35:20]
  wire [7:0] n9_I_34; // @[Top.scala 35:20]
  wire [7:0] n9_I_35; // @[Top.scala 35:20]
  wire [7:0] n9_I_36; // @[Top.scala 35:20]
  wire [7:0] n9_I_37; // @[Top.scala 35:20]
  wire [7:0] n9_I_38; // @[Top.scala 35:20]
  wire [7:0] n9_I_39; // @[Top.scala 35:20]
  wire [7:0] n9_O_0; // @[Top.scala 35:20]
  wire [7:0] n9_O_1; // @[Top.scala 35:20]
  wire [7:0] n9_O_2; // @[Top.scala 35:20]
  wire [7:0] n9_O_3; // @[Top.scala 35:20]
  wire [7:0] n9_O_4; // @[Top.scala 35:20]
  wire [7:0] n9_O_5; // @[Top.scala 35:20]
  wire [7:0] n9_O_6; // @[Top.scala 35:20]
  wire [7:0] n9_O_7; // @[Top.scala 35:20]
  wire [7:0] n9_O_8; // @[Top.scala 35:20]
  wire [7:0] n9_O_9; // @[Top.scala 35:20]
  wire [7:0] n9_O_10; // @[Top.scala 35:20]
  wire [7:0] n9_O_11; // @[Top.scala 35:20]
  wire [7:0] n9_O_12; // @[Top.scala 35:20]
  wire [7:0] n9_O_13; // @[Top.scala 35:20]
  wire [7:0] n9_O_14; // @[Top.scala 35:20]
  wire [7:0] n9_O_15; // @[Top.scala 35:20]
  wire [7:0] n9_O_16; // @[Top.scala 35:20]
  wire [7:0] n9_O_17; // @[Top.scala 35:20]
  wire [7:0] n9_O_18; // @[Top.scala 35:20]
  wire [7:0] n9_O_19; // @[Top.scala 35:20]
  wire [7:0] n9_O_20; // @[Top.scala 35:20]
  wire [7:0] n9_O_21; // @[Top.scala 35:20]
  wire [7:0] n9_O_22; // @[Top.scala 35:20]
  wire [7:0] n9_O_23; // @[Top.scala 35:20]
  wire [7:0] n9_O_24; // @[Top.scala 35:20]
  wire [7:0] n9_O_25; // @[Top.scala 35:20]
  wire [7:0] n9_O_26; // @[Top.scala 35:20]
  wire [7:0] n9_O_27; // @[Top.scala 35:20]
  wire [7:0] n9_O_28; // @[Top.scala 35:20]
  wire [7:0] n9_O_29; // @[Top.scala 35:20]
  wire [7:0] n9_O_30; // @[Top.scala 35:20]
  wire [7:0] n9_O_31; // @[Top.scala 35:20]
  wire [7:0] n9_O_32; // @[Top.scala 35:20]
  wire [7:0] n9_O_33; // @[Top.scala 35:20]
  wire [7:0] n9_O_34; // @[Top.scala 35:20]
  wire [7:0] n9_O_35; // @[Top.scala 35:20]
  wire [7:0] n9_O_36; // @[Top.scala 35:20]
  wire [7:0] n9_O_37; // @[Top.scala 35:20]
  wire [7:0] n9_O_38; // @[Top.scala 35:20]
  wire [7:0] n9_O_39; // @[Top.scala 35:20]
  wire  n10_clock; // @[Top.scala 38:21]
  wire  n10_reset; // @[Top.scala 38:21]
  wire  n10_valid_up; // @[Top.scala 38:21]
  wire  n10_valid_down; // @[Top.scala 38:21]
  wire [7:0] n10_I_0; // @[Top.scala 38:21]
  wire [7:0] n10_I_1; // @[Top.scala 38:21]
  wire [7:0] n10_I_2; // @[Top.scala 38:21]
  wire [7:0] n10_I_3; // @[Top.scala 38:21]
  wire [7:0] n10_I_4; // @[Top.scala 38:21]
  wire [7:0] n10_I_5; // @[Top.scala 38:21]
  wire [7:0] n10_I_6; // @[Top.scala 38:21]
  wire [7:0] n10_I_7; // @[Top.scala 38:21]
  wire [7:0] n10_I_8; // @[Top.scala 38:21]
  wire [7:0] n10_I_9; // @[Top.scala 38:21]
  wire [7:0] n10_I_10; // @[Top.scala 38:21]
  wire [7:0] n10_I_11; // @[Top.scala 38:21]
  wire [7:0] n10_I_12; // @[Top.scala 38:21]
  wire [7:0] n10_I_13; // @[Top.scala 38:21]
  wire [7:0] n10_I_14; // @[Top.scala 38:21]
  wire [7:0] n10_I_15; // @[Top.scala 38:21]
  wire [7:0] n10_I_16; // @[Top.scala 38:21]
  wire [7:0] n10_I_17; // @[Top.scala 38:21]
  wire [7:0] n10_I_18; // @[Top.scala 38:21]
  wire [7:0] n10_I_19; // @[Top.scala 38:21]
  wire [7:0] n10_I_20; // @[Top.scala 38:21]
  wire [7:0] n10_I_21; // @[Top.scala 38:21]
  wire [7:0] n10_I_22; // @[Top.scala 38:21]
  wire [7:0] n10_I_23; // @[Top.scala 38:21]
  wire [7:0] n10_I_24; // @[Top.scala 38:21]
  wire [7:0] n10_I_25; // @[Top.scala 38:21]
  wire [7:0] n10_I_26; // @[Top.scala 38:21]
  wire [7:0] n10_I_27; // @[Top.scala 38:21]
  wire [7:0] n10_I_28; // @[Top.scala 38:21]
  wire [7:0] n10_I_29; // @[Top.scala 38:21]
  wire [7:0] n10_I_30; // @[Top.scala 38:21]
  wire [7:0] n10_I_31; // @[Top.scala 38:21]
  wire [7:0] n10_I_32; // @[Top.scala 38:21]
  wire [7:0] n10_I_33; // @[Top.scala 38:21]
  wire [7:0] n10_I_34; // @[Top.scala 38:21]
  wire [7:0] n10_I_35; // @[Top.scala 38:21]
  wire [7:0] n10_I_36; // @[Top.scala 38:21]
  wire [7:0] n10_I_37; // @[Top.scala 38:21]
  wire [7:0] n10_I_38; // @[Top.scala 38:21]
  wire [7:0] n10_I_39; // @[Top.scala 38:21]
  wire [7:0] n10_O_0; // @[Top.scala 38:21]
  wire [7:0] n10_O_1; // @[Top.scala 38:21]
  wire [7:0] n10_O_2; // @[Top.scala 38:21]
  wire [7:0] n10_O_3; // @[Top.scala 38:21]
  wire [7:0] n10_O_4; // @[Top.scala 38:21]
  wire [7:0] n10_O_5; // @[Top.scala 38:21]
  wire [7:0] n10_O_6; // @[Top.scala 38:21]
  wire [7:0] n10_O_7; // @[Top.scala 38:21]
  wire [7:0] n10_O_8; // @[Top.scala 38:21]
  wire [7:0] n10_O_9; // @[Top.scala 38:21]
  wire [7:0] n10_O_10; // @[Top.scala 38:21]
  wire [7:0] n10_O_11; // @[Top.scala 38:21]
  wire [7:0] n10_O_12; // @[Top.scala 38:21]
  wire [7:0] n10_O_13; // @[Top.scala 38:21]
  wire [7:0] n10_O_14; // @[Top.scala 38:21]
  wire [7:0] n10_O_15; // @[Top.scala 38:21]
  wire [7:0] n10_O_16; // @[Top.scala 38:21]
  wire [7:0] n10_O_17; // @[Top.scala 38:21]
  wire [7:0] n10_O_18; // @[Top.scala 38:21]
  wire [7:0] n10_O_19; // @[Top.scala 38:21]
  wire [7:0] n10_O_20; // @[Top.scala 38:21]
  wire [7:0] n10_O_21; // @[Top.scala 38:21]
  wire [7:0] n10_O_22; // @[Top.scala 38:21]
  wire [7:0] n10_O_23; // @[Top.scala 38:21]
  wire [7:0] n10_O_24; // @[Top.scala 38:21]
  wire [7:0] n10_O_25; // @[Top.scala 38:21]
  wire [7:0] n10_O_26; // @[Top.scala 38:21]
  wire [7:0] n10_O_27; // @[Top.scala 38:21]
  wire [7:0] n10_O_28; // @[Top.scala 38:21]
  wire [7:0] n10_O_29; // @[Top.scala 38:21]
  wire [7:0] n10_O_30; // @[Top.scala 38:21]
  wire [7:0] n10_O_31; // @[Top.scala 38:21]
  wire [7:0] n10_O_32; // @[Top.scala 38:21]
  wire [7:0] n10_O_33; // @[Top.scala 38:21]
  wire [7:0] n10_O_34; // @[Top.scala 38:21]
  wire [7:0] n10_O_35; // @[Top.scala 38:21]
  wire [7:0] n10_O_36; // @[Top.scala 38:21]
  wire [7:0] n10_O_37; // @[Top.scala 38:21]
  wire [7:0] n10_O_38; // @[Top.scala 38:21]
  wire [7:0] n10_O_39; // @[Top.scala 38:21]
  wire  n11_clock; // @[Top.scala 41:21]
  wire  n11_reset; // @[Top.scala 41:21]
  wire  n11_valid_up; // @[Top.scala 41:21]
  wire  n11_valid_down; // @[Top.scala 41:21]
  wire [7:0] n11_I_0; // @[Top.scala 41:21]
  wire [7:0] n11_I_1; // @[Top.scala 41:21]
  wire [7:0] n11_I_2; // @[Top.scala 41:21]
  wire [7:0] n11_I_3; // @[Top.scala 41:21]
  wire [7:0] n11_I_4; // @[Top.scala 41:21]
  wire [7:0] n11_I_5; // @[Top.scala 41:21]
  wire [7:0] n11_I_6; // @[Top.scala 41:21]
  wire [7:0] n11_I_7; // @[Top.scala 41:21]
  wire [7:0] n11_I_8; // @[Top.scala 41:21]
  wire [7:0] n11_I_9; // @[Top.scala 41:21]
  wire [7:0] n11_I_10; // @[Top.scala 41:21]
  wire [7:0] n11_I_11; // @[Top.scala 41:21]
  wire [7:0] n11_I_12; // @[Top.scala 41:21]
  wire [7:0] n11_I_13; // @[Top.scala 41:21]
  wire [7:0] n11_I_14; // @[Top.scala 41:21]
  wire [7:0] n11_I_15; // @[Top.scala 41:21]
  wire [7:0] n11_I_16; // @[Top.scala 41:21]
  wire [7:0] n11_I_17; // @[Top.scala 41:21]
  wire [7:0] n11_I_18; // @[Top.scala 41:21]
  wire [7:0] n11_I_19; // @[Top.scala 41:21]
  wire [7:0] n11_I_20; // @[Top.scala 41:21]
  wire [7:0] n11_I_21; // @[Top.scala 41:21]
  wire [7:0] n11_I_22; // @[Top.scala 41:21]
  wire [7:0] n11_I_23; // @[Top.scala 41:21]
  wire [7:0] n11_I_24; // @[Top.scala 41:21]
  wire [7:0] n11_I_25; // @[Top.scala 41:21]
  wire [7:0] n11_I_26; // @[Top.scala 41:21]
  wire [7:0] n11_I_27; // @[Top.scala 41:21]
  wire [7:0] n11_I_28; // @[Top.scala 41:21]
  wire [7:0] n11_I_29; // @[Top.scala 41:21]
  wire [7:0] n11_I_30; // @[Top.scala 41:21]
  wire [7:0] n11_I_31; // @[Top.scala 41:21]
  wire [7:0] n11_I_32; // @[Top.scala 41:21]
  wire [7:0] n11_I_33; // @[Top.scala 41:21]
  wire [7:0] n11_I_34; // @[Top.scala 41:21]
  wire [7:0] n11_I_35; // @[Top.scala 41:21]
  wire [7:0] n11_I_36; // @[Top.scala 41:21]
  wire [7:0] n11_I_37; // @[Top.scala 41:21]
  wire [7:0] n11_I_38; // @[Top.scala 41:21]
  wire [7:0] n11_I_39; // @[Top.scala 41:21]
  wire [7:0] n11_O_0; // @[Top.scala 41:21]
  wire [7:0] n11_O_1; // @[Top.scala 41:21]
  wire [7:0] n11_O_2; // @[Top.scala 41:21]
  wire [7:0] n11_O_3; // @[Top.scala 41:21]
  wire [7:0] n11_O_4; // @[Top.scala 41:21]
  wire [7:0] n11_O_5; // @[Top.scala 41:21]
  wire [7:0] n11_O_6; // @[Top.scala 41:21]
  wire [7:0] n11_O_7; // @[Top.scala 41:21]
  wire [7:0] n11_O_8; // @[Top.scala 41:21]
  wire [7:0] n11_O_9; // @[Top.scala 41:21]
  wire [7:0] n11_O_10; // @[Top.scala 41:21]
  wire [7:0] n11_O_11; // @[Top.scala 41:21]
  wire [7:0] n11_O_12; // @[Top.scala 41:21]
  wire [7:0] n11_O_13; // @[Top.scala 41:21]
  wire [7:0] n11_O_14; // @[Top.scala 41:21]
  wire [7:0] n11_O_15; // @[Top.scala 41:21]
  wire [7:0] n11_O_16; // @[Top.scala 41:21]
  wire [7:0] n11_O_17; // @[Top.scala 41:21]
  wire [7:0] n11_O_18; // @[Top.scala 41:21]
  wire [7:0] n11_O_19; // @[Top.scala 41:21]
  wire [7:0] n11_O_20; // @[Top.scala 41:21]
  wire [7:0] n11_O_21; // @[Top.scala 41:21]
  wire [7:0] n11_O_22; // @[Top.scala 41:21]
  wire [7:0] n11_O_23; // @[Top.scala 41:21]
  wire [7:0] n11_O_24; // @[Top.scala 41:21]
  wire [7:0] n11_O_25; // @[Top.scala 41:21]
  wire [7:0] n11_O_26; // @[Top.scala 41:21]
  wire [7:0] n11_O_27; // @[Top.scala 41:21]
  wire [7:0] n11_O_28; // @[Top.scala 41:21]
  wire [7:0] n11_O_29; // @[Top.scala 41:21]
  wire [7:0] n11_O_30; // @[Top.scala 41:21]
  wire [7:0] n11_O_31; // @[Top.scala 41:21]
  wire [7:0] n11_O_32; // @[Top.scala 41:21]
  wire [7:0] n11_O_33; // @[Top.scala 41:21]
  wire [7:0] n11_O_34; // @[Top.scala 41:21]
  wire [7:0] n11_O_35; // @[Top.scala 41:21]
  wire [7:0] n11_O_36; // @[Top.scala 41:21]
  wire [7:0] n11_O_37; // @[Top.scala 41:21]
  wire [7:0] n11_O_38; // @[Top.scala 41:21]
  wire [7:0] n11_O_39; // @[Top.scala 41:21]
  wire  n12_clock; // @[Top.scala 44:21]
  wire  n12_reset; // @[Top.scala 44:21]
  wire  n12_valid_up; // @[Top.scala 44:21]
  wire  n12_valid_down; // @[Top.scala 44:21]
  wire [7:0] n12_I_0; // @[Top.scala 44:21]
  wire [7:0] n12_I_1; // @[Top.scala 44:21]
  wire [7:0] n12_I_2; // @[Top.scala 44:21]
  wire [7:0] n12_I_3; // @[Top.scala 44:21]
  wire [7:0] n12_I_4; // @[Top.scala 44:21]
  wire [7:0] n12_I_5; // @[Top.scala 44:21]
  wire [7:0] n12_I_6; // @[Top.scala 44:21]
  wire [7:0] n12_I_7; // @[Top.scala 44:21]
  wire [7:0] n12_I_8; // @[Top.scala 44:21]
  wire [7:0] n12_I_9; // @[Top.scala 44:21]
  wire [7:0] n12_I_10; // @[Top.scala 44:21]
  wire [7:0] n12_I_11; // @[Top.scala 44:21]
  wire [7:0] n12_I_12; // @[Top.scala 44:21]
  wire [7:0] n12_I_13; // @[Top.scala 44:21]
  wire [7:0] n12_I_14; // @[Top.scala 44:21]
  wire [7:0] n12_I_15; // @[Top.scala 44:21]
  wire [7:0] n12_I_16; // @[Top.scala 44:21]
  wire [7:0] n12_I_17; // @[Top.scala 44:21]
  wire [7:0] n12_I_18; // @[Top.scala 44:21]
  wire [7:0] n12_I_19; // @[Top.scala 44:21]
  wire [7:0] n12_I_20; // @[Top.scala 44:21]
  wire [7:0] n12_I_21; // @[Top.scala 44:21]
  wire [7:0] n12_I_22; // @[Top.scala 44:21]
  wire [7:0] n12_I_23; // @[Top.scala 44:21]
  wire [7:0] n12_I_24; // @[Top.scala 44:21]
  wire [7:0] n12_I_25; // @[Top.scala 44:21]
  wire [7:0] n12_I_26; // @[Top.scala 44:21]
  wire [7:0] n12_I_27; // @[Top.scala 44:21]
  wire [7:0] n12_I_28; // @[Top.scala 44:21]
  wire [7:0] n12_I_29; // @[Top.scala 44:21]
  wire [7:0] n12_I_30; // @[Top.scala 44:21]
  wire [7:0] n12_I_31; // @[Top.scala 44:21]
  wire [7:0] n12_I_32; // @[Top.scala 44:21]
  wire [7:0] n12_I_33; // @[Top.scala 44:21]
  wire [7:0] n12_I_34; // @[Top.scala 44:21]
  wire [7:0] n12_I_35; // @[Top.scala 44:21]
  wire [7:0] n12_I_36; // @[Top.scala 44:21]
  wire [7:0] n12_I_37; // @[Top.scala 44:21]
  wire [7:0] n12_I_38; // @[Top.scala 44:21]
  wire [7:0] n12_I_39; // @[Top.scala 44:21]
  wire [7:0] n12_O_0; // @[Top.scala 44:21]
  wire [7:0] n12_O_1; // @[Top.scala 44:21]
  wire [7:0] n12_O_2; // @[Top.scala 44:21]
  wire [7:0] n12_O_3; // @[Top.scala 44:21]
  wire [7:0] n12_O_4; // @[Top.scala 44:21]
  wire [7:0] n12_O_5; // @[Top.scala 44:21]
  wire [7:0] n12_O_6; // @[Top.scala 44:21]
  wire [7:0] n12_O_7; // @[Top.scala 44:21]
  wire [7:0] n12_O_8; // @[Top.scala 44:21]
  wire [7:0] n12_O_9; // @[Top.scala 44:21]
  wire [7:0] n12_O_10; // @[Top.scala 44:21]
  wire [7:0] n12_O_11; // @[Top.scala 44:21]
  wire [7:0] n12_O_12; // @[Top.scala 44:21]
  wire [7:0] n12_O_13; // @[Top.scala 44:21]
  wire [7:0] n12_O_14; // @[Top.scala 44:21]
  wire [7:0] n12_O_15; // @[Top.scala 44:21]
  wire [7:0] n12_O_16; // @[Top.scala 44:21]
  wire [7:0] n12_O_17; // @[Top.scala 44:21]
  wire [7:0] n12_O_18; // @[Top.scala 44:21]
  wire [7:0] n12_O_19; // @[Top.scala 44:21]
  wire [7:0] n12_O_20; // @[Top.scala 44:21]
  wire [7:0] n12_O_21; // @[Top.scala 44:21]
  wire [7:0] n12_O_22; // @[Top.scala 44:21]
  wire [7:0] n12_O_23; // @[Top.scala 44:21]
  wire [7:0] n12_O_24; // @[Top.scala 44:21]
  wire [7:0] n12_O_25; // @[Top.scala 44:21]
  wire [7:0] n12_O_26; // @[Top.scala 44:21]
  wire [7:0] n12_O_27; // @[Top.scala 44:21]
  wire [7:0] n12_O_28; // @[Top.scala 44:21]
  wire [7:0] n12_O_29; // @[Top.scala 44:21]
  wire [7:0] n12_O_30; // @[Top.scala 44:21]
  wire [7:0] n12_O_31; // @[Top.scala 44:21]
  wire [7:0] n12_O_32; // @[Top.scala 44:21]
  wire [7:0] n12_O_33; // @[Top.scala 44:21]
  wire [7:0] n12_O_34; // @[Top.scala 44:21]
  wire [7:0] n12_O_35; // @[Top.scala 44:21]
  wire [7:0] n12_O_36; // @[Top.scala 44:21]
  wire [7:0] n12_O_37; // @[Top.scala 44:21]
  wire [7:0] n12_O_38; // @[Top.scala 44:21]
  wire [7:0] n12_O_39; // @[Top.scala 44:21]
  FIFO n1 ( // @[Top.scala 32:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .I_8(n1_I_8),
    .I_9(n1_I_9),
    .I_10(n1_I_10),
    .I_11(n1_I_11),
    .I_12(n1_I_12),
    .I_13(n1_I_13),
    .I_14(n1_I_14),
    .I_15(n1_I_15),
    .I_16(n1_I_16),
    .I_17(n1_I_17),
    .I_18(n1_I_18),
    .I_19(n1_I_19),
    .I_20(n1_I_20),
    .I_21(n1_I_21),
    .I_22(n1_I_22),
    .I_23(n1_I_23),
    .I_24(n1_I_24),
    .I_25(n1_I_25),
    .I_26(n1_I_26),
    .I_27(n1_I_27),
    .I_28(n1_I_28),
    .I_29(n1_I_29),
    .I_30(n1_I_30),
    .I_31(n1_I_31),
    .I_32(n1_I_32),
    .I_33(n1_I_33),
    .I_34(n1_I_34),
    .I_35(n1_I_35),
    .I_36(n1_I_36),
    .I_37(n1_I_37),
    .I_38(n1_I_38),
    .I_39(n1_I_39),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7),
    .O_8(n1_O_8),
    .O_9(n1_O_9),
    .O_10(n1_O_10),
    .O_11(n1_O_11),
    .O_12(n1_O_12),
    .O_13(n1_O_13),
    .O_14(n1_O_14),
    .O_15(n1_O_15),
    .O_16(n1_O_16),
    .O_17(n1_O_17),
    .O_18(n1_O_18),
    .O_19(n1_O_19),
    .O_20(n1_O_20),
    .O_21(n1_O_21),
    .O_22(n1_O_22),
    .O_23(n1_O_23),
    .O_24(n1_O_24),
    .O_25(n1_O_25),
    .O_26(n1_O_26),
    .O_27(n1_O_27),
    .O_28(n1_O_28),
    .O_29(n1_O_29),
    .O_30(n1_O_30),
    .O_31(n1_O_31),
    .O_32(n1_O_32),
    .O_33(n1_O_33),
    .O_34(n1_O_34),
    .O_35(n1_O_35),
    .O_36(n1_O_36),
    .O_37(n1_O_37),
    .O_38(n1_O_38),
    .O_39(n1_O_39)
  );
  MapT n9 ( // @[Top.scala 35:20]
    .clock(n9_clock),
    .reset(n9_reset),
    .valid_up(n9_valid_up),
    .valid_down(n9_valid_down),
    .I_0(n9_I_0),
    .I_1(n9_I_1),
    .I_2(n9_I_2),
    .I_3(n9_I_3),
    .I_4(n9_I_4),
    .I_5(n9_I_5),
    .I_6(n9_I_6),
    .I_7(n9_I_7),
    .I_8(n9_I_8),
    .I_9(n9_I_9),
    .I_10(n9_I_10),
    .I_11(n9_I_11),
    .I_12(n9_I_12),
    .I_13(n9_I_13),
    .I_14(n9_I_14),
    .I_15(n9_I_15),
    .I_16(n9_I_16),
    .I_17(n9_I_17),
    .I_18(n9_I_18),
    .I_19(n9_I_19),
    .I_20(n9_I_20),
    .I_21(n9_I_21),
    .I_22(n9_I_22),
    .I_23(n9_I_23),
    .I_24(n9_I_24),
    .I_25(n9_I_25),
    .I_26(n9_I_26),
    .I_27(n9_I_27),
    .I_28(n9_I_28),
    .I_29(n9_I_29),
    .I_30(n9_I_30),
    .I_31(n9_I_31),
    .I_32(n9_I_32),
    .I_33(n9_I_33),
    .I_34(n9_I_34),
    .I_35(n9_I_35),
    .I_36(n9_I_36),
    .I_37(n9_I_37),
    .I_38(n9_I_38),
    .I_39(n9_I_39),
    .O_0(n9_O_0),
    .O_1(n9_O_1),
    .O_2(n9_O_2),
    .O_3(n9_O_3),
    .O_4(n9_O_4),
    .O_5(n9_O_5),
    .O_6(n9_O_6),
    .O_7(n9_O_7),
    .O_8(n9_O_8),
    .O_9(n9_O_9),
    .O_10(n9_O_10),
    .O_11(n9_O_11),
    .O_12(n9_O_12),
    .O_13(n9_O_13),
    .O_14(n9_O_14),
    .O_15(n9_O_15),
    .O_16(n9_O_16),
    .O_17(n9_O_17),
    .O_18(n9_O_18),
    .O_19(n9_O_19),
    .O_20(n9_O_20),
    .O_21(n9_O_21),
    .O_22(n9_O_22),
    .O_23(n9_O_23),
    .O_24(n9_O_24),
    .O_25(n9_O_25),
    .O_26(n9_O_26),
    .O_27(n9_O_27),
    .O_28(n9_O_28),
    .O_29(n9_O_29),
    .O_30(n9_O_30),
    .O_31(n9_O_31),
    .O_32(n9_O_32),
    .O_33(n9_O_33),
    .O_34(n9_O_34),
    .O_35(n9_O_35),
    .O_36(n9_O_36),
    .O_37(n9_O_37),
    .O_38(n9_O_38),
    .O_39(n9_O_39)
  );
  FIFO n10 ( // @[Top.scala 38:21]
    .clock(n10_clock),
    .reset(n10_reset),
    .valid_up(n10_valid_up),
    .valid_down(n10_valid_down),
    .I_0(n10_I_0),
    .I_1(n10_I_1),
    .I_2(n10_I_2),
    .I_3(n10_I_3),
    .I_4(n10_I_4),
    .I_5(n10_I_5),
    .I_6(n10_I_6),
    .I_7(n10_I_7),
    .I_8(n10_I_8),
    .I_9(n10_I_9),
    .I_10(n10_I_10),
    .I_11(n10_I_11),
    .I_12(n10_I_12),
    .I_13(n10_I_13),
    .I_14(n10_I_14),
    .I_15(n10_I_15),
    .I_16(n10_I_16),
    .I_17(n10_I_17),
    .I_18(n10_I_18),
    .I_19(n10_I_19),
    .I_20(n10_I_20),
    .I_21(n10_I_21),
    .I_22(n10_I_22),
    .I_23(n10_I_23),
    .I_24(n10_I_24),
    .I_25(n10_I_25),
    .I_26(n10_I_26),
    .I_27(n10_I_27),
    .I_28(n10_I_28),
    .I_29(n10_I_29),
    .I_30(n10_I_30),
    .I_31(n10_I_31),
    .I_32(n10_I_32),
    .I_33(n10_I_33),
    .I_34(n10_I_34),
    .I_35(n10_I_35),
    .I_36(n10_I_36),
    .I_37(n10_I_37),
    .I_38(n10_I_38),
    .I_39(n10_I_39),
    .O_0(n10_O_0),
    .O_1(n10_O_1),
    .O_2(n10_O_2),
    .O_3(n10_O_3),
    .O_4(n10_O_4),
    .O_5(n10_O_5),
    .O_6(n10_O_6),
    .O_7(n10_O_7),
    .O_8(n10_O_8),
    .O_9(n10_O_9),
    .O_10(n10_O_10),
    .O_11(n10_O_11),
    .O_12(n10_O_12),
    .O_13(n10_O_13),
    .O_14(n10_O_14),
    .O_15(n10_O_15),
    .O_16(n10_O_16),
    .O_17(n10_O_17),
    .O_18(n10_O_18),
    .O_19(n10_O_19),
    .O_20(n10_O_20),
    .O_21(n10_O_21),
    .O_22(n10_O_22),
    .O_23(n10_O_23),
    .O_24(n10_O_24),
    .O_25(n10_O_25),
    .O_26(n10_O_26),
    .O_27(n10_O_27),
    .O_28(n10_O_28),
    .O_29(n10_O_29),
    .O_30(n10_O_30),
    .O_31(n10_O_31),
    .O_32(n10_O_32),
    .O_33(n10_O_33),
    .O_34(n10_O_34),
    .O_35(n10_O_35),
    .O_36(n10_O_36),
    .O_37(n10_O_37),
    .O_38(n10_O_38),
    .O_39(n10_O_39)
  );
  FIFO n11 ( // @[Top.scala 41:21]
    .clock(n11_clock),
    .reset(n11_reset),
    .valid_up(n11_valid_up),
    .valid_down(n11_valid_down),
    .I_0(n11_I_0),
    .I_1(n11_I_1),
    .I_2(n11_I_2),
    .I_3(n11_I_3),
    .I_4(n11_I_4),
    .I_5(n11_I_5),
    .I_6(n11_I_6),
    .I_7(n11_I_7),
    .I_8(n11_I_8),
    .I_9(n11_I_9),
    .I_10(n11_I_10),
    .I_11(n11_I_11),
    .I_12(n11_I_12),
    .I_13(n11_I_13),
    .I_14(n11_I_14),
    .I_15(n11_I_15),
    .I_16(n11_I_16),
    .I_17(n11_I_17),
    .I_18(n11_I_18),
    .I_19(n11_I_19),
    .I_20(n11_I_20),
    .I_21(n11_I_21),
    .I_22(n11_I_22),
    .I_23(n11_I_23),
    .I_24(n11_I_24),
    .I_25(n11_I_25),
    .I_26(n11_I_26),
    .I_27(n11_I_27),
    .I_28(n11_I_28),
    .I_29(n11_I_29),
    .I_30(n11_I_30),
    .I_31(n11_I_31),
    .I_32(n11_I_32),
    .I_33(n11_I_33),
    .I_34(n11_I_34),
    .I_35(n11_I_35),
    .I_36(n11_I_36),
    .I_37(n11_I_37),
    .I_38(n11_I_38),
    .I_39(n11_I_39),
    .O_0(n11_O_0),
    .O_1(n11_O_1),
    .O_2(n11_O_2),
    .O_3(n11_O_3),
    .O_4(n11_O_4),
    .O_5(n11_O_5),
    .O_6(n11_O_6),
    .O_7(n11_O_7),
    .O_8(n11_O_8),
    .O_9(n11_O_9),
    .O_10(n11_O_10),
    .O_11(n11_O_11),
    .O_12(n11_O_12),
    .O_13(n11_O_13),
    .O_14(n11_O_14),
    .O_15(n11_O_15),
    .O_16(n11_O_16),
    .O_17(n11_O_17),
    .O_18(n11_O_18),
    .O_19(n11_O_19),
    .O_20(n11_O_20),
    .O_21(n11_O_21),
    .O_22(n11_O_22),
    .O_23(n11_O_23),
    .O_24(n11_O_24),
    .O_25(n11_O_25),
    .O_26(n11_O_26),
    .O_27(n11_O_27),
    .O_28(n11_O_28),
    .O_29(n11_O_29),
    .O_30(n11_O_30),
    .O_31(n11_O_31),
    .O_32(n11_O_32),
    .O_33(n11_O_33),
    .O_34(n11_O_34),
    .O_35(n11_O_35),
    .O_36(n11_O_36),
    .O_37(n11_O_37),
    .O_38(n11_O_38),
    .O_39(n11_O_39)
  );
  FIFO n12 ( // @[Top.scala 44:21]
    .clock(n12_clock),
    .reset(n12_reset),
    .valid_up(n12_valid_up),
    .valid_down(n12_valid_down),
    .I_0(n12_I_0),
    .I_1(n12_I_1),
    .I_2(n12_I_2),
    .I_3(n12_I_3),
    .I_4(n12_I_4),
    .I_5(n12_I_5),
    .I_6(n12_I_6),
    .I_7(n12_I_7),
    .I_8(n12_I_8),
    .I_9(n12_I_9),
    .I_10(n12_I_10),
    .I_11(n12_I_11),
    .I_12(n12_I_12),
    .I_13(n12_I_13),
    .I_14(n12_I_14),
    .I_15(n12_I_15),
    .I_16(n12_I_16),
    .I_17(n12_I_17),
    .I_18(n12_I_18),
    .I_19(n12_I_19),
    .I_20(n12_I_20),
    .I_21(n12_I_21),
    .I_22(n12_I_22),
    .I_23(n12_I_23),
    .I_24(n12_I_24),
    .I_25(n12_I_25),
    .I_26(n12_I_26),
    .I_27(n12_I_27),
    .I_28(n12_I_28),
    .I_29(n12_I_29),
    .I_30(n12_I_30),
    .I_31(n12_I_31),
    .I_32(n12_I_32),
    .I_33(n12_I_33),
    .I_34(n12_I_34),
    .I_35(n12_I_35),
    .I_36(n12_I_36),
    .I_37(n12_I_37),
    .I_38(n12_I_38),
    .I_39(n12_I_39),
    .O_0(n12_O_0),
    .O_1(n12_O_1),
    .O_2(n12_O_2),
    .O_3(n12_O_3),
    .O_4(n12_O_4),
    .O_5(n12_O_5),
    .O_6(n12_O_6),
    .O_7(n12_O_7),
    .O_8(n12_O_8),
    .O_9(n12_O_9),
    .O_10(n12_O_10),
    .O_11(n12_O_11),
    .O_12(n12_O_12),
    .O_13(n12_O_13),
    .O_14(n12_O_14),
    .O_15(n12_O_15),
    .O_16(n12_O_16),
    .O_17(n12_O_17),
    .O_18(n12_O_18),
    .O_19(n12_O_19),
    .O_20(n12_O_20),
    .O_21(n12_O_21),
    .O_22(n12_O_22),
    .O_23(n12_O_23),
    .O_24(n12_O_24),
    .O_25(n12_O_25),
    .O_26(n12_O_26),
    .O_27(n12_O_27),
    .O_28(n12_O_28),
    .O_29(n12_O_29),
    .O_30(n12_O_30),
    .O_31(n12_O_31),
    .O_32(n12_O_32),
    .O_33(n12_O_33),
    .O_34(n12_O_34),
    .O_35(n12_O_35),
    .O_36(n12_O_36),
    .O_37(n12_O_37),
    .O_38(n12_O_38),
    .O_39(n12_O_39)
  );
  assign valid_down = n12_valid_down; // @[Top.scala 48:16]
  assign O_0 = n12_O_0; // @[Top.scala 47:7]
  assign O_1 = n12_O_1; // @[Top.scala 47:7]
  assign O_2 = n12_O_2; // @[Top.scala 47:7]
  assign O_3 = n12_O_3; // @[Top.scala 47:7]
  assign O_4 = n12_O_4; // @[Top.scala 47:7]
  assign O_5 = n12_O_5; // @[Top.scala 47:7]
  assign O_6 = n12_O_6; // @[Top.scala 47:7]
  assign O_7 = n12_O_7; // @[Top.scala 47:7]
  assign O_8 = n12_O_8; // @[Top.scala 47:7]
  assign O_9 = n12_O_9; // @[Top.scala 47:7]
  assign O_10 = n12_O_10; // @[Top.scala 47:7]
  assign O_11 = n12_O_11; // @[Top.scala 47:7]
  assign O_12 = n12_O_12; // @[Top.scala 47:7]
  assign O_13 = n12_O_13; // @[Top.scala 47:7]
  assign O_14 = n12_O_14; // @[Top.scala 47:7]
  assign O_15 = n12_O_15; // @[Top.scala 47:7]
  assign O_16 = n12_O_16; // @[Top.scala 47:7]
  assign O_17 = n12_O_17; // @[Top.scala 47:7]
  assign O_18 = n12_O_18; // @[Top.scala 47:7]
  assign O_19 = n12_O_19; // @[Top.scala 47:7]
  assign O_20 = n12_O_20; // @[Top.scala 47:7]
  assign O_21 = n12_O_21; // @[Top.scala 47:7]
  assign O_22 = n12_O_22; // @[Top.scala 47:7]
  assign O_23 = n12_O_23; // @[Top.scala 47:7]
  assign O_24 = n12_O_24; // @[Top.scala 47:7]
  assign O_25 = n12_O_25; // @[Top.scala 47:7]
  assign O_26 = n12_O_26; // @[Top.scala 47:7]
  assign O_27 = n12_O_27; // @[Top.scala 47:7]
  assign O_28 = n12_O_28; // @[Top.scala 47:7]
  assign O_29 = n12_O_29; // @[Top.scala 47:7]
  assign O_30 = n12_O_30; // @[Top.scala 47:7]
  assign O_31 = n12_O_31; // @[Top.scala 47:7]
  assign O_32 = n12_O_32; // @[Top.scala 47:7]
  assign O_33 = n12_O_33; // @[Top.scala 47:7]
  assign O_34 = n12_O_34; // @[Top.scala 47:7]
  assign O_35 = n12_O_35; // @[Top.scala 47:7]
  assign O_36 = n12_O_36; // @[Top.scala 47:7]
  assign O_37 = n12_O_37; // @[Top.scala 47:7]
  assign O_38 = n12_O_38; // @[Top.scala 47:7]
  assign O_39 = n12_O_39; // @[Top.scala 47:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 34:17]
  assign n1_I_0 = I_0; // @[Top.scala 33:10]
  assign n1_I_1 = I_1; // @[Top.scala 33:10]
  assign n1_I_2 = I_2; // @[Top.scala 33:10]
  assign n1_I_3 = I_3; // @[Top.scala 33:10]
  assign n1_I_4 = I_4; // @[Top.scala 33:10]
  assign n1_I_5 = I_5; // @[Top.scala 33:10]
  assign n1_I_6 = I_6; // @[Top.scala 33:10]
  assign n1_I_7 = I_7; // @[Top.scala 33:10]
  assign n1_I_8 = I_8; // @[Top.scala 33:10]
  assign n1_I_9 = I_9; // @[Top.scala 33:10]
  assign n1_I_10 = I_10; // @[Top.scala 33:10]
  assign n1_I_11 = I_11; // @[Top.scala 33:10]
  assign n1_I_12 = I_12; // @[Top.scala 33:10]
  assign n1_I_13 = I_13; // @[Top.scala 33:10]
  assign n1_I_14 = I_14; // @[Top.scala 33:10]
  assign n1_I_15 = I_15; // @[Top.scala 33:10]
  assign n1_I_16 = I_16; // @[Top.scala 33:10]
  assign n1_I_17 = I_17; // @[Top.scala 33:10]
  assign n1_I_18 = I_18; // @[Top.scala 33:10]
  assign n1_I_19 = I_19; // @[Top.scala 33:10]
  assign n1_I_20 = I_20; // @[Top.scala 33:10]
  assign n1_I_21 = I_21; // @[Top.scala 33:10]
  assign n1_I_22 = I_22; // @[Top.scala 33:10]
  assign n1_I_23 = I_23; // @[Top.scala 33:10]
  assign n1_I_24 = I_24; // @[Top.scala 33:10]
  assign n1_I_25 = I_25; // @[Top.scala 33:10]
  assign n1_I_26 = I_26; // @[Top.scala 33:10]
  assign n1_I_27 = I_27; // @[Top.scala 33:10]
  assign n1_I_28 = I_28; // @[Top.scala 33:10]
  assign n1_I_29 = I_29; // @[Top.scala 33:10]
  assign n1_I_30 = I_30; // @[Top.scala 33:10]
  assign n1_I_31 = I_31; // @[Top.scala 33:10]
  assign n1_I_32 = I_32; // @[Top.scala 33:10]
  assign n1_I_33 = I_33; // @[Top.scala 33:10]
  assign n1_I_34 = I_34; // @[Top.scala 33:10]
  assign n1_I_35 = I_35; // @[Top.scala 33:10]
  assign n1_I_36 = I_36; // @[Top.scala 33:10]
  assign n1_I_37 = I_37; // @[Top.scala 33:10]
  assign n1_I_38 = I_38; // @[Top.scala 33:10]
  assign n1_I_39 = I_39; // @[Top.scala 33:10]
  assign n9_clock = clock;
  assign n9_reset = reset;
  assign n9_valid_up = n1_valid_down; // @[Top.scala 37:17]
  assign n9_I_0 = n1_O_0; // @[Top.scala 36:10]
  assign n9_I_1 = n1_O_1; // @[Top.scala 36:10]
  assign n9_I_2 = n1_O_2; // @[Top.scala 36:10]
  assign n9_I_3 = n1_O_3; // @[Top.scala 36:10]
  assign n9_I_4 = n1_O_4; // @[Top.scala 36:10]
  assign n9_I_5 = n1_O_5; // @[Top.scala 36:10]
  assign n9_I_6 = n1_O_6; // @[Top.scala 36:10]
  assign n9_I_7 = n1_O_7; // @[Top.scala 36:10]
  assign n9_I_8 = n1_O_8; // @[Top.scala 36:10]
  assign n9_I_9 = n1_O_9; // @[Top.scala 36:10]
  assign n9_I_10 = n1_O_10; // @[Top.scala 36:10]
  assign n9_I_11 = n1_O_11; // @[Top.scala 36:10]
  assign n9_I_12 = n1_O_12; // @[Top.scala 36:10]
  assign n9_I_13 = n1_O_13; // @[Top.scala 36:10]
  assign n9_I_14 = n1_O_14; // @[Top.scala 36:10]
  assign n9_I_15 = n1_O_15; // @[Top.scala 36:10]
  assign n9_I_16 = n1_O_16; // @[Top.scala 36:10]
  assign n9_I_17 = n1_O_17; // @[Top.scala 36:10]
  assign n9_I_18 = n1_O_18; // @[Top.scala 36:10]
  assign n9_I_19 = n1_O_19; // @[Top.scala 36:10]
  assign n9_I_20 = n1_O_20; // @[Top.scala 36:10]
  assign n9_I_21 = n1_O_21; // @[Top.scala 36:10]
  assign n9_I_22 = n1_O_22; // @[Top.scala 36:10]
  assign n9_I_23 = n1_O_23; // @[Top.scala 36:10]
  assign n9_I_24 = n1_O_24; // @[Top.scala 36:10]
  assign n9_I_25 = n1_O_25; // @[Top.scala 36:10]
  assign n9_I_26 = n1_O_26; // @[Top.scala 36:10]
  assign n9_I_27 = n1_O_27; // @[Top.scala 36:10]
  assign n9_I_28 = n1_O_28; // @[Top.scala 36:10]
  assign n9_I_29 = n1_O_29; // @[Top.scala 36:10]
  assign n9_I_30 = n1_O_30; // @[Top.scala 36:10]
  assign n9_I_31 = n1_O_31; // @[Top.scala 36:10]
  assign n9_I_32 = n1_O_32; // @[Top.scala 36:10]
  assign n9_I_33 = n1_O_33; // @[Top.scala 36:10]
  assign n9_I_34 = n1_O_34; // @[Top.scala 36:10]
  assign n9_I_35 = n1_O_35; // @[Top.scala 36:10]
  assign n9_I_36 = n1_O_36; // @[Top.scala 36:10]
  assign n9_I_37 = n1_O_37; // @[Top.scala 36:10]
  assign n9_I_38 = n1_O_38; // @[Top.scala 36:10]
  assign n9_I_39 = n1_O_39; // @[Top.scala 36:10]
  assign n10_clock = clock;
  assign n10_reset = reset;
  assign n10_valid_up = n9_valid_down; // @[Top.scala 40:18]
  assign n10_I_0 = n9_O_0; // @[Top.scala 39:11]
  assign n10_I_1 = n9_O_1; // @[Top.scala 39:11]
  assign n10_I_2 = n9_O_2; // @[Top.scala 39:11]
  assign n10_I_3 = n9_O_3; // @[Top.scala 39:11]
  assign n10_I_4 = n9_O_4; // @[Top.scala 39:11]
  assign n10_I_5 = n9_O_5; // @[Top.scala 39:11]
  assign n10_I_6 = n9_O_6; // @[Top.scala 39:11]
  assign n10_I_7 = n9_O_7; // @[Top.scala 39:11]
  assign n10_I_8 = n9_O_8; // @[Top.scala 39:11]
  assign n10_I_9 = n9_O_9; // @[Top.scala 39:11]
  assign n10_I_10 = n9_O_10; // @[Top.scala 39:11]
  assign n10_I_11 = n9_O_11; // @[Top.scala 39:11]
  assign n10_I_12 = n9_O_12; // @[Top.scala 39:11]
  assign n10_I_13 = n9_O_13; // @[Top.scala 39:11]
  assign n10_I_14 = n9_O_14; // @[Top.scala 39:11]
  assign n10_I_15 = n9_O_15; // @[Top.scala 39:11]
  assign n10_I_16 = n9_O_16; // @[Top.scala 39:11]
  assign n10_I_17 = n9_O_17; // @[Top.scala 39:11]
  assign n10_I_18 = n9_O_18; // @[Top.scala 39:11]
  assign n10_I_19 = n9_O_19; // @[Top.scala 39:11]
  assign n10_I_20 = n9_O_20; // @[Top.scala 39:11]
  assign n10_I_21 = n9_O_21; // @[Top.scala 39:11]
  assign n10_I_22 = n9_O_22; // @[Top.scala 39:11]
  assign n10_I_23 = n9_O_23; // @[Top.scala 39:11]
  assign n10_I_24 = n9_O_24; // @[Top.scala 39:11]
  assign n10_I_25 = n9_O_25; // @[Top.scala 39:11]
  assign n10_I_26 = n9_O_26; // @[Top.scala 39:11]
  assign n10_I_27 = n9_O_27; // @[Top.scala 39:11]
  assign n10_I_28 = n9_O_28; // @[Top.scala 39:11]
  assign n10_I_29 = n9_O_29; // @[Top.scala 39:11]
  assign n10_I_30 = n9_O_30; // @[Top.scala 39:11]
  assign n10_I_31 = n9_O_31; // @[Top.scala 39:11]
  assign n10_I_32 = n9_O_32; // @[Top.scala 39:11]
  assign n10_I_33 = n9_O_33; // @[Top.scala 39:11]
  assign n10_I_34 = n9_O_34; // @[Top.scala 39:11]
  assign n10_I_35 = n9_O_35; // @[Top.scala 39:11]
  assign n10_I_36 = n9_O_36; // @[Top.scala 39:11]
  assign n10_I_37 = n9_O_37; // @[Top.scala 39:11]
  assign n10_I_38 = n9_O_38; // @[Top.scala 39:11]
  assign n10_I_39 = n9_O_39; // @[Top.scala 39:11]
  assign n11_clock = clock;
  assign n11_reset = reset;
  assign n11_valid_up = n10_valid_down; // @[Top.scala 43:18]
  assign n11_I_0 = n10_O_0; // @[Top.scala 42:11]
  assign n11_I_1 = n10_O_1; // @[Top.scala 42:11]
  assign n11_I_2 = n10_O_2; // @[Top.scala 42:11]
  assign n11_I_3 = n10_O_3; // @[Top.scala 42:11]
  assign n11_I_4 = n10_O_4; // @[Top.scala 42:11]
  assign n11_I_5 = n10_O_5; // @[Top.scala 42:11]
  assign n11_I_6 = n10_O_6; // @[Top.scala 42:11]
  assign n11_I_7 = n10_O_7; // @[Top.scala 42:11]
  assign n11_I_8 = n10_O_8; // @[Top.scala 42:11]
  assign n11_I_9 = n10_O_9; // @[Top.scala 42:11]
  assign n11_I_10 = n10_O_10; // @[Top.scala 42:11]
  assign n11_I_11 = n10_O_11; // @[Top.scala 42:11]
  assign n11_I_12 = n10_O_12; // @[Top.scala 42:11]
  assign n11_I_13 = n10_O_13; // @[Top.scala 42:11]
  assign n11_I_14 = n10_O_14; // @[Top.scala 42:11]
  assign n11_I_15 = n10_O_15; // @[Top.scala 42:11]
  assign n11_I_16 = n10_O_16; // @[Top.scala 42:11]
  assign n11_I_17 = n10_O_17; // @[Top.scala 42:11]
  assign n11_I_18 = n10_O_18; // @[Top.scala 42:11]
  assign n11_I_19 = n10_O_19; // @[Top.scala 42:11]
  assign n11_I_20 = n10_O_20; // @[Top.scala 42:11]
  assign n11_I_21 = n10_O_21; // @[Top.scala 42:11]
  assign n11_I_22 = n10_O_22; // @[Top.scala 42:11]
  assign n11_I_23 = n10_O_23; // @[Top.scala 42:11]
  assign n11_I_24 = n10_O_24; // @[Top.scala 42:11]
  assign n11_I_25 = n10_O_25; // @[Top.scala 42:11]
  assign n11_I_26 = n10_O_26; // @[Top.scala 42:11]
  assign n11_I_27 = n10_O_27; // @[Top.scala 42:11]
  assign n11_I_28 = n10_O_28; // @[Top.scala 42:11]
  assign n11_I_29 = n10_O_29; // @[Top.scala 42:11]
  assign n11_I_30 = n10_O_30; // @[Top.scala 42:11]
  assign n11_I_31 = n10_O_31; // @[Top.scala 42:11]
  assign n11_I_32 = n10_O_32; // @[Top.scala 42:11]
  assign n11_I_33 = n10_O_33; // @[Top.scala 42:11]
  assign n11_I_34 = n10_O_34; // @[Top.scala 42:11]
  assign n11_I_35 = n10_O_35; // @[Top.scala 42:11]
  assign n11_I_36 = n10_O_36; // @[Top.scala 42:11]
  assign n11_I_37 = n10_O_37; // @[Top.scala 42:11]
  assign n11_I_38 = n10_O_38; // @[Top.scala 42:11]
  assign n11_I_39 = n10_O_39; // @[Top.scala 42:11]
  assign n12_clock = clock;
  assign n12_reset = reset;
  assign n12_valid_up = n11_valid_down; // @[Top.scala 46:18]
  assign n12_I_0 = n11_O_0; // @[Top.scala 45:11]
  assign n12_I_1 = n11_O_1; // @[Top.scala 45:11]
  assign n12_I_2 = n11_O_2; // @[Top.scala 45:11]
  assign n12_I_3 = n11_O_3; // @[Top.scala 45:11]
  assign n12_I_4 = n11_O_4; // @[Top.scala 45:11]
  assign n12_I_5 = n11_O_5; // @[Top.scala 45:11]
  assign n12_I_6 = n11_O_6; // @[Top.scala 45:11]
  assign n12_I_7 = n11_O_7; // @[Top.scala 45:11]
  assign n12_I_8 = n11_O_8; // @[Top.scala 45:11]
  assign n12_I_9 = n11_O_9; // @[Top.scala 45:11]
  assign n12_I_10 = n11_O_10; // @[Top.scala 45:11]
  assign n12_I_11 = n11_O_11; // @[Top.scala 45:11]
  assign n12_I_12 = n11_O_12; // @[Top.scala 45:11]
  assign n12_I_13 = n11_O_13; // @[Top.scala 45:11]
  assign n12_I_14 = n11_O_14; // @[Top.scala 45:11]
  assign n12_I_15 = n11_O_15; // @[Top.scala 45:11]
  assign n12_I_16 = n11_O_16; // @[Top.scala 45:11]
  assign n12_I_17 = n11_O_17; // @[Top.scala 45:11]
  assign n12_I_18 = n11_O_18; // @[Top.scala 45:11]
  assign n12_I_19 = n11_O_19; // @[Top.scala 45:11]
  assign n12_I_20 = n11_O_20; // @[Top.scala 45:11]
  assign n12_I_21 = n11_O_21; // @[Top.scala 45:11]
  assign n12_I_22 = n11_O_22; // @[Top.scala 45:11]
  assign n12_I_23 = n11_O_23; // @[Top.scala 45:11]
  assign n12_I_24 = n11_O_24; // @[Top.scala 45:11]
  assign n12_I_25 = n11_O_25; // @[Top.scala 45:11]
  assign n12_I_26 = n11_O_26; // @[Top.scala 45:11]
  assign n12_I_27 = n11_O_27; // @[Top.scala 45:11]
  assign n12_I_28 = n11_O_28; // @[Top.scala 45:11]
  assign n12_I_29 = n11_O_29; // @[Top.scala 45:11]
  assign n12_I_30 = n11_O_30; // @[Top.scala 45:11]
  assign n12_I_31 = n11_O_31; // @[Top.scala 45:11]
  assign n12_I_32 = n11_O_32; // @[Top.scala 45:11]
  assign n12_I_33 = n11_O_33; // @[Top.scala 45:11]
  assign n12_I_34 = n11_O_34; // @[Top.scala 45:11]
  assign n12_I_35 = n11_O_35; // @[Top.scala 45:11]
  assign n12_I_36 = n11_O_36; // @[Top.scala 45:11]
  assign n12_I_37 = n11_O_37; // @[Top.scala 45:11]
  assign n12_I_38 = n11_O_38; // @[Top.scala 45:11]
  assign n12_I_39 = n11_O_39; // @[Top.scala 45:11]
endmodule
