module corebit_and (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 & in1;
endmodule

module atomTupleCreator_t0Int_t1Int (input [7:0] I0/*verilator public*/, input [7:0] I1/*verilator public*/, output [7:0] O__0/*verilator public*/, output [7:0] O__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O__0 = I0;
assign O__1 = I1;
assign valid_down = valid_up;
endmodule

module coreir_ult #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 < in1;
endmodule

module coreir_term #(parameter width = 1) (input [width-1:0] in/*verilator public*/);

endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk/*verilator public*/, input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  reg [width-1:0] outReg/*verilator public*/=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_mux #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, input sel/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = sel ? in1 : in0;
endmodule

module coreir_eq #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 == in1;
endmodule

module coreir_const #(parameter width = 1, parameter value = 1) (output [width-1:0] out/*verilator public*/);
  assign out = value;
endmodule

module coreir_add #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = in0 + in1;
endmodule

module \commonlib_muxn__N2__width1 (input [0:0] in_data_0/*verilator public*/, input [0:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [0:0] out/*verilator public*/);
wire [0:0] _join_out;
coreir_mux #(.width(1)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module lutN #(parameter N = 1, parameter init = 1) (input [N-1:0] in/*verilator public*/, output out/*verilator public*/);
  assign out = init[in];
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit8 (input [7:0] in/*verilator public*/, output [7:0] out/*verilator public*/);
assign out = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit (input in/*verilator public*/, output [0:0] out/*verilator public*/);
assign out = in;
endmodule

module Term_Bitt (input I/*verilator public*/);
wire [0:0] dehydrate_tBit_inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
coreir_term #(.width(1)) term_w1_inst0(.in(dehydrate_tBit_inst0_out));
endmodule

module SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/);
wire [0:0] const_0_1_out;
Term_Bitt Term_Bitt_inst0(.I(CE));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
assign O = const_0_1_out;
endmodule

module Mux2xOutBits1 (input [0:0] I0/*verilator public*/, input [0:0] I1/*verilator public*/, output [0:0] O/*verilator public*/, input S/*verilator public*/);
wire [0:0] coreir_commonlib_mux2x1_inst0_out;
\commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x1_inst0_out));
assign O = coreir_commonlib_mux2x1_inst0_out;
endmodule

module Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1 (input CE/*verilator public*/, input CLK/*verilator public*/, input [0:0] I/*verilator public*/, output [0:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [0:0] Mux2xOutBits1_inst0_O;
wire [0:0] const_0_1_out;
wire [0:0] enable_mux_O;
wire [0:0] value_out;
Mux2xOutBits1 Mux2xOutBits1_inst0(.I0(enable_mux_O), .I1(const_0_1_out), .O(Mux2xOutBits1_inst0_O), .S(RESET));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
Mux2xOutBits1 enable_mux(.I0(value_out), .I1(I), .O(enable_mux_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) value(.clk(CLK), .in(Mux2xOutBits1_inst0_O), .out(value_out));
assign O = value_out;
endmodule

module LUT1_2 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h2), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_1 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h1), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_0 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h0), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT_Array_8_Bit_t_1n (input CLK/*verilator public*/, input [0:0] addr/*verilator public*/, output [7:0] data/*verilator public*/);
wire LUT1_0_inst0_O;
wire LUT1_0_inst1_O;
wire LUT1_0_inst2_O;
wire LUT1_0_inst3_O;
wire LUT1_0_inst4_O;
wire LUT1_0_inst5_O;
wire LUT1_1_inst0_O;
wire LUT1_1_inst1_O;
wire [7:0] hydrate_tArray_8_Bit__inst0_out;
LUT1_0 LUT1_0_inst0(.I0(addr[0]), .O(LUT1_0_inst0_O));
LUT1_0 LUT1_0_inst1(.I0(addr[0]), .O(LUT1_0_inst1_O));
LUT1_0 LUT1_0_inst2(.I0(addr[0]), .O(LUT1_0_inst2_O));
LUT1_0 LUT1_0_inst3(.I0(addr[0]), .O(LUT1_0_inst3_O));
LUT1_0 LUT1_0_inst4(.I0(addr[0]), .O(LUT1_0_inst4_O));
LUT1_0 LUT1_0_inst5(.I0(addr[0]), .O(LUT1_0_inst5_O));
LUT1_1 LUT1_1_inst0(.I0(addr[0]), .O(LUT1_1_inst0_O));
LUT1_1 LUT1_1_inst1(.I0(addr[0]), .O(LUT1_1_inst1_O));
\aetherlinglib_hydrate__hydratedTypeBit8 hydrate_tArray_8_Bit__inst0(.in({LUT1_0_inst5_O,LUT1_0_inst4_O,LUT1_0_inst3_O,LUT1_0_inst2_O,LUT1_0_inst1_O,LUT1_1_inst1_O,LUT1_0_inst0_O,LUT1_1_inst0_O}), .out(hydrate_tArray_8_Bit__inst0_out));
assign data = hydrate_tArray_8_Bit__inst0_out;
endmodule

module DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Register8 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_8_Bit_t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] Register8_inst0_O;
Register8 Register8_inst0(.CLK(CLK), .I(I), .O(Register8_inst0_O));
assign O = Register8_inst0_O;
endmodule

module Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/);
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9_O;
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(I_0), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1(.CLK(CLK), .I(I_1), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10(.CLK(CLK), .I(I_10), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11(.CLK(CLK), .I(I_11), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12(.CLK(CLK), .I(I_12), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13(.CLK(CLK), .I(I_13), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14(.CLK(CLK), .I(I_14), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15(.CLK(CLK), .I(I_15), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16(.CLK(CLK), .I(I_16), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17(.CLK(CLK), .I(I_17), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18(.CLK(CLK), .I(I_18), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19(.CLK(CLK), .I(I_19), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2(.CLK(CLK), .I(I_2), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3(.CLK(CLK), .I(I_3), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4(.CLK(CLK), .I(I_4), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5(.CLK(CLK), .I(I_5), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6(.CLK(CLK), .I(I_6), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7(.CLK(CLK), .I(I_7), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8(.CLK(CLK), .I(I_8), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9(.CLK(CLK), .I(I_9), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9_O));
assign O_0 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
assign O_1 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O;
assign O_10 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10_O;
assign O_11 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11_O;
assign O_12 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12_O;
assign O_13 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13_O;
assign O_14 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14_O;
assign O_15 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15_O;
assign O_16 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16_O;
assign O_17 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17_O;
assign O_18 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18_O;
assign O_19 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19_O;
assign O_2 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O;
assign O_3 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3_O;
assign O_4 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4_O;
assign O_5 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5_O;
assign O_6 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6_O;
assign O_7 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7_O;
assign O_8 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8_O;
assign O_9 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9_O;
endmodule

module Register1 (input CLK/*verilator public*/, input [0:0] I/*verilator public*/, output [0:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
assign O = DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
endmodule

module Register_Bitt_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] Register1_inst0_O;
Register1 Register1_inst0(.CLK(CLK), .I(I), .O(Register1_inst0_O));
assign O = Register1_inst0_O[0];
endmodule

module FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
wire [7:0] Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_11(I_11), .I_12(I_12), .I_13(I_13), .I_14(I_14), .I_15(I_15), .I_16(I_16), .I_17(I_17), .I_18(I_18), .I_19(I_19), .I_2(I_2), .I_3(I_3), .I_4(I_4), .I_5(I_5), .I_6(I_6), .I_7(I_7), .I_8(I_8), .I_9(I_9), .O_0(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0), .O_1(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1), .O_10(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10), .O_11(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11), .O_12(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12), .O_13(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13), .O_14(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14), .O_15(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15), .O_16(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16), .O_17(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17), .O_18(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18), .O_19(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19), .O_2(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2), .O_3(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3), .O_4(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4), .O_5(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5), .O_6(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6), .O_7(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7), .O_8(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8), .O_9(Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign O_1 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
assign O_10 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
assign O_11 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
assign O_12 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
assign O_13 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
assign O_14 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
assign O_15 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
assign O_16 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
assign O_17 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
assign O_18 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
assign O_19 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
assign O_2 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
assign O_3 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
assign O_4 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
assign O_5 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
assign O_6 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
assign O_7 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
assign O_8 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
assign O_9 = Register_Array_20_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Counter1CER (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [0:0] Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O;
wire [0:0] const_1_1_out;
wire [0:0] coreir_add1_inst0_out;
Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1 Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0(.CE(CE), .CLK(CLK), .I(coreir_add1_inst0_out), .O(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O), .RESET(RESET));
coreir_const #(.value(1'h1), .width(1)) const_1_1(.out(const_1_1_out));
coreir_add #(.width(1)) coreir_add1_inst0(.in0(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O), .in1(const_1_1_out), .out(coreir_add1_inst0_out));
assign O = Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O;
endmodule

module Counter1_Mod2CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/);
wire [0:0] Counter1CER_inst0_O;
wire LUT1_2_inst0_O;
wire and_inst0_out;
Counter1CER Counter1CER_inst0(.CE(CE), .CLK(CLK), .O(Counter1CER_inst0_O), .RESET(and_inst0_out));
LUT1_2 LUT1_2_inst0(.I0(Counter1CER_inst0_O[0]), .O(LUT1_2_inst0_O));
corebit_and and_inst0(.in0(LUT1_2_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter1CER_inst0_O;
endmodule

module InitialDelayCounter_1 (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [0:0] Counter1_Mod2CE_inst0_O;
wire and_inst0_out;
wire [0:0] coreir_const11_inst0_out;
wire coreir_eq_1_inst0_out;
wire coreir_ult1_inst0_out;
Counter1_Mod2CE Counter1_Mod2CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter1_Mod2CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult1_inst0_out), .out(and_inst0_out));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
coreir_eq #(.width(1)) coreir_eq_1_inst0(.in0(Counter1_Mod2CE_inst0_O), .in1(coreir_const11_inst0_out), .out(coreir_eq_1_inst0_out));
coreir_ult #(.width(1)) coreir_ult1_inst0(.in0(Counter1_Mod2CE_inst0_O), .in1(coreir_const11_inst0_out), .out(coreir_ult1_inst0_out));
assign valid = coreir_eq_1_inst0_out;
endmodule

module Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire InitialDelayCounter_1_inst0_valid;
wire [7:0] LUT_Array_8_Bit_t_1n_inst0_data;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
InitialDelayCounter_1 InitialDelayCounter_1_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_1_inst0_valid));
LUT_Array_8_Bit_t_1n LUT_Array_8_Bit_t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data(LUT_Array_8_Bit_t_1n_inst0_data));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(InitialDelayCounter_1_inst0_valid), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O = LUT_Array_8_Bit_t_1n_inst0_data;
assign valid_down = InitialDelayCounter_1_inst0_valid;
endmodule

module Add_Atom (input [7:0] I__0/*verilator public*/, input [7:0] I__1/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] coreir_add8_inst0_out;
coreir_add #(.width(8)) coreir_add8_inst0(.in0(I__0), .in1(I__1), .out(coreir_add8_inst0_out));
assign O = coreir_add8_inst0_out;
assign valid_down = valid_up;
endmodule

module Module_0 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Add_Atom_inst0_O;
wire Add_Atom_inst0_valid_down;
wire [7:0] Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O;
wire Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire and_inst0_out;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
Add_Atom Add_Atom_inst0(.I__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .I__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .O(Add_Atom_inst0_O), .valid_down(Add_Atom_inst0_valid_down), .valid_up(atomTupleCreator_t0Int_t1Int_inst0_valid_down));
Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .valid_down(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(valid_up), .in1(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I), .I1(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(and_inst0_out));
assign O = Add_Atom_inst0_O;
assign valid_down = Add_Atom_inst0_valid_down;
endmodule

module NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Module_0_inst0_O;
wire Module_0_inst0_valid_down;
wire [7:0] Module_0_inst1_O;
wire Module_0_inst1_valid_down;
wire [7:0] Module_0_inst10_O;
wire Module_0_inst10_valid_down;
wire [7:0] Module_0_inst11_O;
wire Module_0_inst11_valid_down;
wire [7:0] Module_0_inst12_O;
wire Module_0_inst12_valid_down;
wire [7:0] Module_0_inst13_O;
wire Module_0_inst13_valid_down;
wire [7:0] Module_0_inst14_O;
wire Module_0_inst14_valid_down;
wire [7:0] Module_0_inst15_O;
wire Module_0_inst15_valid_down;
wire [7:0] Module_0_inst16_O;
wire Module_0_inst16_valid_down;
wire [7:0] Module_0_inst17_O;
wire Module_0_inst17_valid_down;
wire [7:0] Module_0_inst18_O;
wire Module_0_inst18_valid_down;
wire [7:0] Module_0_inst19_O;
wire Module_0_inst19_valid_down;
wire [7:0] Module_0_inst2_O;
wire Module_0_inst2_valid_down;
wire [7:0] Module_0_inst3_O;
wire Module_0_inst3_valid_down;
wire [7:0] Module_0_inst4_O;
wire Module_0_inst4_valid_down;
wire [7:0] Module_0_inst5_O;
wire Module_0_inst5_valid_down;
wire [7:0] Module_0_inst6_O;
wire Module_0_inst6_valid_down;
wire [7:0] Module_0_inst7_O;
wire Module_0_inst7_valid_down;
wire [7:0] Module_0_inst8_O;
wire Module_0_inst8_valid_down;
wire [7:0] Module_0_inst9_O;
wire Module_0_inst9_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst11_out;
wire and_inst12_out;
wire and_inst13_out;
wire and_inst14_out;
wire and_inst15_out;
wire and_inst16_out;
wire and_inst17_out;
wire and_inst18_out;
wire and_inst2_out;
wire and_inst3_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
wire and_inst8_out;
wire and_inst9_out;
Module_0 Module_0_inst0(.CLK(CLK), .I(I_0), .O(Module_0_inst0_O), .valid_down(Module_0_inst0_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst1(.CLK(CLK), .I(I_1), .O(Module_0_inst1_O), .valid_down(Module_0_inst1_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst10(.CLK(CLK), .I(I_10), .O(Module_0_inst10_O), .valid_down(Module_0_inst10_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst11(.CLK(CLK), .I(I_11), .O(Module_0_inst11_O), .valid_down(Module_0_inst11_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst12(.CLK(CLK), .I(I_12), .O(Module_0_inst12_O), .valid_down(Module_0_inst12_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst13(.CLK(CLK), .I(I_13), .O(Module_0_inst13_O), .valid_down(Module_0_inst13_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst14(.CLK(CLK), .I(I_14), .O(Module_0_inst14_O), .valid_down(Module_0_inst14_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst15(.CLK(CLK), .I(I_15), .O(Module_0_inst15_O), .valid_down(Module_0_inst15_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst16(.CLK(CLK), .I(I_16), .O(Module_0_inst16_O), .valid_down(Module_0_inst16_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst17(.CLK(CLK), .I(I_17), .O(Module_0_inst17_O), .valid_down(Module_0_inst17_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst18(.CLK(CLK), .I(I_18), .O(Module_0_inst18_O), .valid_down(Module_0_inst18_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst19(.CLK(CLK), .I(I_19), .O(Module_0_inst19_O), .valid_down(Module_0_inst19_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst2(.CLK(CLK), .I(I_2), .O(Module_0_inst2_O), .valid_down(Module_0_inst2_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst3(.CLK(CLK), .I(I_3), .O(Module_0_inst3_O), .valid_down(Module_0_inst3_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst4(.CLK(CLK), .I(I_4), .O(Module_0_inst4_O), .valid_down(Module_0_inst4_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst5(.CLK(CLK), .I(I_5), .O(Module_0_inst5_O), .valid_down(Module_0_inst5_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst6(.CLK(CLK), .I(I_6), .O(Module_0_inst6_O), .valid_down(Module_0_inst6_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst7(.CLK(CLK), .I(I_7), .O(Module_0_inst7_O), .valid_down(Module_0_inst7_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst8(.CLK(CLK), .I(I_8), .O(Module_0_inst8_O), .valid_down(Module_0_inst8_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst9(.CLK(CLK), .I(I_9), .O(Module_0_inst9_O), .valid_down(Module_0_inst9_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Module_0_inst0_valid_down), .in1(Module_0_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Module_0_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(Module_0_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(Module_0_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(Module_0_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(Module_0_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(Module_0_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(Module_0_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(Module_0_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(Module_0_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(Module_0_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Module_0_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Module_0_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Module_0_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Module_0_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Module_0_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Module_0_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(Module_0_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(Module_0_inst10_valid_down), .out(and_inst9_out));
assign O_0 = Module_0_inst0_O;
assign O_1 = Module_0_inst1_O;
assign O_10 = Module_0_inst10_O;
assign O_11 = Module_0_inst11_O;
assign O_12 = Module_0_inst12_O;
assign O_13 = Module_0_inst13_O;
assign O_14 = Module_0_inst14_O;
assign O_15 = Module_0_inst15_O;
assign O_16 = Module_0_inst16_O;
assign O_17 = Module_0_inst17_O;
assign O_18 = Module_0_inst18_O;
assign O_19 = Module_0_inst19_O;
assign O_2 = Module_0_inst2_O;
assign O_3 = Module_0_inst3_O;
assign O_4 = Module_0_inst4_O;
assign O_5 = Module_0_inst5_O;
assign O_6 = Module_0_inst6_O;
assign O_7 = Module_0_inst7_O;
assign O_8 = Module_0_inst8_O;
assign O_9 = Module_0_inst9_O;
assign valid_down = and_inst18_out;
endmodule

module Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
wire [7:0] NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
wire NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_11(I_11), .I_12(I_12), .I_13(I_13), .I_14(I_14), .I_15(I_15), .I_16(I_16), .I_17(I_17), .I_18(I_18), .I_19(I_19), .I_2(I_2), .I_3(I_3), .I_4(I_4), .I_5(I_5), .I_6(I_6), .I_7(I_7), .I_8(I_8), .I_9(I_9), .O_0(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_10(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .O_11(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .O_12(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .O_13(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .O_14(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .O_15(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .O_16(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .O_17(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .O_18(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .O_19(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .O_2(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .O_3(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .O_4(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .O_5(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .O_6(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .O_7(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .O_8(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .O_9(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .valid_down(NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
assign O_1 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
assign O_10 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
assign O_11 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
assign O_12 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
assign O_13 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
assign O_14 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
assign O_15 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
assign O_16 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
assign O_17 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
assign O_18 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
assign O_19 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
assign O_2 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
assign O_3 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
assign O_4 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
assign O_5 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
assign O_6 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
assign O_7 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
assign O_8 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
assign O_9 = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
assign valid_down = NativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module top (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9;
wire FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9;
wire FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9;
wire FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9;
wire FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_0;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_1;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_10;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_11;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_12;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_13;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_14;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_15;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_16;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_17;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_18;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_19;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_2;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_3;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_4;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_5;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_6;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_7;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_8;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_9;
wire FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_valid_down;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_0;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_1;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_10;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_11;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_12;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_13;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_14;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_15;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_16;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_17;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_18;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_19;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_2;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_3;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_4;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_5;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_6;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_7;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_8;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_9;
wire FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_valid_down;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_0;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_1;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_10;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_11;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_12;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_13;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_14;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_15;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_16;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_17;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_18;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_19;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_2;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_3;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_4;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_5;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_6;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_7;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_8;
wire [7:0] FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_9;
wire FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_valid_down;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
wire [7:0] Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
wire Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_11(I_11), .I_12(I_12), .I_13(I_13), .I_14(I_14), .I_15(I_15), .I_16(I_16), .I_17(I_17), .I_18(I_18), .I_19(I_19), .I_2(I_2), .I_3(I_3), .I_4(I_4), .I_5(I_5), .I_6(I_6), .I_7(I_7), .I_8(I_8), .I_9(I_9), .O_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .O_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .O_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .O_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .O_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .O_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .O_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .O_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .O_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .O_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .O_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .O_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .O_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .O_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .O_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .O_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .O_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .valid_down(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .I_1(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .I_10(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .I_11(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .I_12(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .I_13(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .I_14(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .I_15(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .I_16(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .I_17(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .I_18(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .I_19(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .I_2(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .I_3(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .I_4(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .I_5(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .I_6(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .I_7(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .I_8(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .I_9(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .O_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .O_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .O_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .O_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .O_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .O_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .O_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .O_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .O_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .O_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .O_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .O_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .O_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .O_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .O_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .O_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .O_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .O_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .O_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .O_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .valid_down(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down));
FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .I_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .I_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .I_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .I_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .I_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .I_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .I_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .I_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .I_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .I_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .I_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .I_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .I_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .I_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .I_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .I_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .I_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .I_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .I_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .O_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1), .O_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10), .O_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11), .O_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12), .O_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13), .O_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14), .O_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15), .O_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16), .O_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17), .O_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18), .O_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19), .O_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2), .O_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3), .O_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4), .O_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5), .O_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6), .O_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7), .O_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8), .O_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9), .valid_down(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down));
FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3(.CLK(CLK), .I_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .I_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1), .I_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10), .I_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11), .I_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12), .I_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13), .I_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14), .I_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15), .I_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16), .I_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17), .I_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18), .I_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19), .I_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2), .I_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3), .I_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4), .I_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5), .I_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6), .I_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7), .I_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8), .I_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9), .O_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .O_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1), .O_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10), .O_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11), .O_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12), .O_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13), .O_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14), .O_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15), .O_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16), .O_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17), .O_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18), .O_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19), .O_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2), .O_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3), .O_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4), .O_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5), .O_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6), .O_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7), .O_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8), .O_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9), .valid_down(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down), .valid_up(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down));
FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4(.CLK(CLK), .I_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .I_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1), .I_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10), .I_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11), .I_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12), .I_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13), .I_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14), .I_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15), .I_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16), .I_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17), .I_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18), .I_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19), .I_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2), .I_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3), .I_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4), .I_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5), .I_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6), .I_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7), .I_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8), .I_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9), .O_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_0), .O_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_1), .O_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_10), .O_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_11), .O_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_12), .O_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_13), .O_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_14), .O_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_15), .O_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_16), .O_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_17), .O_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_18), .O_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_19), .O_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_2), .O_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_3), .O_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_4), .O_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_5), .O_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_6), .O_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_7), .O_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_8), .O_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_9), .valid_down(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_valid_down), .valid_up(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down));
FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5(.CLK(CLK), .I_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_0), .I_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_1), .I_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_10), .I_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_11), .I_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_12), .I_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_13), .I_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_14), .I_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_15), .I_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_16), .I_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_17), .I_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_18), .I_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_19), .I_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_2), .I_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_3), .I_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_4), .I_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_5), .I_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_6), .I_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_7), .I_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_8), .I_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_O_9), .O_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_0), .O_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_1), .O_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_10), .O_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_11), .O_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_12), .O_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_13), .O_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_14), .O_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_15), .O_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_16), .O_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_17), .O_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_18), .O_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_19), .O_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_2), .O_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_3), .O_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_4), .O_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_5), .O_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_6), .O_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_7), .O_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_8), .O_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_9), .valid_down(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_valid_down), .valid_up(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst4_valid_down));
FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6(.CLK(CLK), .I_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_0), .I_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_1), .I_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_10), .I_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_11), .I_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_12), .I_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_13), .I_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_14), .I_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_15), .I_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_16), .I_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_17), .I_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_18), .I_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_19), .I_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_2), .I_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_3), .I_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_4), .I_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_5), .I_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_6), .I_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_7), .I_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_8), .I_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_O_9), .O_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_0), .O_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_1), .O_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_10), .O_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_11), .O_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_12), .O_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_13), .O_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_14), .O_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_15), .O_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_16), .O_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_17), .O_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_18), .O_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_19), .O_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_2), .O_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_3), .O_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_4), .O_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_5), .O_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_6), .O_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_7), .O_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_8), .O_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_9), .valid_down(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_valid_down), .valid_up(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst5_valid_down));
Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0(.CLK(CLK), .I_0(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I_1(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I_10(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .I_11(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .I_12(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .I_13(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .I_14(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .I_15(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .I_16(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .I_17(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .I_18(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .I_19(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .I_2(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .I_3(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .I_4(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .I_5(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .I_6(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .I_7(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .I_8(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .I_9(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .O_0(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_10(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .O_11(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .O_12(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .O_13(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .O_14(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .O_15(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .O_16(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .O_17(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .O_18(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .O_19(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .O_2(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .O_3(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .O_4(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .O_5(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .O_6(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .O_7(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .O_8(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .O_9(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .valid_down(Map_T_n10_i0_opNativeMapParallel_n20_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_20_Array_8_In_Bit____O_Array_20_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
assign O_0 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_0;
assign O_1 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_1;
assign O_10 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_10;
assign O_11 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_11;
assign O_12 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_12;
assign O_13 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_13;
assign O_14 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_14;
assign O_15 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_15;
assign O_16 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_16;
assign O_17 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_17;
assign O_18 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_18;
assign O_19 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_19;
assign O_2 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_2;
assign O_3 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_3;
assign O_4 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_4;
assign O_5 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_5;
assign O_6 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_6;
assign O_7 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_7;
assign O_8 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_8;
assign O_9 = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_O_9;
assign valid_down = FIFO_tTSeq_10_0_SSeq_20_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst6_valid_down;
endmodule

